--CPLD oR FPGA
--WS2812BCLK .=. 0.4us
--WS2812B�X�ʾ�

Library IEEE;						--�s���s��w
Use IEEE.std_logic_1164.all;		--�ޥήM��
Use IEEE.std_logic_unsigned.all;	--�ޥήM��

entity WS2812B_Driver is
	port(	WS2812BCLK,WS2812BRESET,loadck:in std_logic;--�ާ@�W�v,���m,���Jck
			LEDGRBdata:in std_logic_vector(23 downto 0);--��m���
			reload,emitter,WS2812Bout:out std_logic		--�n�D���J,�o�g���A,�o�g��X 
		);
end entity WS2812B_Driver;

architecture Albert of WS2812B_Driver is
	signal load_clr,reload1:std_logic:='0';	--���J�H���ާ@
	signal LEDGRBdata0,LEDGRBdata1:std_logic_vector(23 downto 0);--��m��Ƹ��J
	signal DATA01:std_logic_vector(2 downto 0):="000";			 --�s�X�줸:bit out=>0:100,1:110
	signal DATAn:integer range 0 to 31:=0;	--��m��Ʀ줸����
	signal bitn:integer range 0 to 3:=0;	--�s�X�줸�o�g��

begin

WS2812Bout<=DATA01(2);--LED��m��Ʀ줸��X
reload<=not (reload1 or load_clr) and WS2812BRESET;--�w�ľ��n�D���J��Ư߽�

--�w���w�ľ�--------------------
LEDdata_load:
process(loadck,WS2812BRESET)
begin
	if WS2812BRESET='0' or (load_clr='1' and reload1='1') then
		reload1<='0'; --�w�ľ���
	elsif rising_edge(loadck) then	--��m��Ƹ��Jck
		LEDGRBdata1<=LEDGRBdata;	--��m��Ƹ��J�w�ľ�
		reload1<='1';--�w�ľ���
	end if;		
end process LEDdata_load;

WS2812B_Send:process(WS2812BCLK,WS2812BRESET)
begin
	if WS2812BRESET='0' then
		DATA01<="000";	--��X����줸
		load_clr<='0';	--���\�w�ľ��ʧ@
		emitter<='0';	--����o�g
		DATAn<=0;		--���ݵo�g�줸��
		bitn<=0;		--�s�X�줸�o�g��0�줸
	elsif rising_edge(WS2812BCLK) then
		load_clr<='0';						--���\�w�ľ��ʧ@
		if bitn/=0 then			--�|���s�X�줸���o�g
			DATA01<=DATA01(1 downto 0) & "0";--�o�g�줸
			bitn<=bitn-1;					 --�s�X�줸�o�g�줸��1
		elsif DATAn/=0 then		--�|����Ʀ줸���s�X
			DATA01<='1' & LEDGRBdata0(DATAn-1) & '0';--�o�g�줸�s�X(���ݵo�g�줸�s�X��3�줸)
			DATAn<=DATAn-1;				--���ݵo�g�줸�ƴ�1
			bitn<=2;					--�s�X�줸�o�g��2�줸
		elsif reload1='1' then	--�w�ľ��w����m��ƶi��
			LEDGRBdata0<=LEDGRBdata1;	--��m��Ƹ��J
			DATAn<=23;					--���ݵo�g�줸��
			DATA01<='1' & LEDGRBdata1(23) & '0';--�o�g�줸�s�X(���ݵo�g�줸�s�X��3�줸)
			bitn<=2;					--�s�X�줸�o�g��2�줸
			load_clr<='1';				--�w���J�o�g��,�M���w�ľ�
			emitter<='1';				--�o�g��
		else					--�w�ľ��L��m���
			emitter<='0';				--����o�g
		end if;
	end if;
end process WS2812B_Send;

end Albert;
