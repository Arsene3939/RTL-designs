--MG90S ����
--EP3C16Q240C8 50MHz LEs:15,408 PINs:161 ,gckp31 ,SResetp99

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;


entity MG90S_Driver is
	port(MG90S_CLK,MG90S_RESET:in std_logic;	--MG90S_Driver�X��clk(6.25MHz),reset�H��
		 MG90S_dir0:in std_logic;				--��ʤ�V0
		 MG90S_deg0:in integer range 0 to 90;	--��ʨ���0
		 MG90S_o0:out std_logic;				--Driver��X1
		 MG90S_dir1:in std_logic;				--��ʤ�V1
		 MG90S_deg1:in integer range 0 to 90;	--��ʨ���1
		 MG90S_o1:out std_logic);				--Driver��X1
end MG90S_Driver;

architecture Albert of MG90S_Driver is
	signal MG90Servo:integer range 0 to 125000;	--servo pwm���;�
	
	--MG90Servopwm ���(function(��'0'�t'1',��0~90)) 
	function MG90Servopwm(MG90S_dir:in std_logic;MG90S_deg:in integer range 0 to 90) return integer is
		variable MG90Servod:integer range 0 to 6000;--3125; --���״����
		variable MG90Servos:integer range 0 to 16000;--12500;--servo pwm��v��
		begin
			--MG90Servod:=347*MG90S_deg/10;	--���״����
			
			MG90Servod:=380*MG90S_deg/6;	--���״����(�g�ץ���)
			if MG90S_dir='0' then
				MG90Servos:=9375+MG90Servod;--servo pwm��v��
			else
				MG90Servos:=9375-MG90Servod;--servo pwm��v��
			end if;
			return MG90Servos;
	end MG90Servopwm;

-- --------------------------
begin
--servo pwm���;�--------------------------------------------------
MG90S_o0<='1' when MG90Servo<MG90Servopwm(MG90S_dir0,MG90S_deg0) and MG90S_RESET='1' else '0';
MG90S_o1<='1' when MG90Servo<MG90Servopwm(MG90S_dir1,MG90S_deg1) and MG90S_RESET='1' else '0';
MG90S:process(MG90S_CLK,MG90S_RESET)
begin
	if MG90S_RESET='0' then
		MG90Servo<=0;
	elsif rising_edge(MG90S_CLK) then
		MG90Servo<=MG90Servo+1;
		if MG90Servo=124999 then
			MG90Servo<=0;
		end if;
	end if;
end Process MG90S;

end Albert;
