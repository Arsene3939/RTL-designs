--Dht11_Driver
--Data format:
--DHT11_DBo(std_logic_vector:8bit):��DHT11_RDp�����X��
--RDp=5:chK_SUM
--RDp=4							   3							   2								1								  0					
--The 8bit humidity integer data + 8bit the Humidity decimal data +8 bit temperature integer data + 8bit fractional temperature data +8 bit parity bit.
--������X���(DHT11_DBoH)�ηū�(DHT11_DBoT):integer(0~255:8bit)
--107.01.01��
--EP3C16Q240C8 50MHz

Library IEEE;						--�s���s��w
Use IEEE.std_logic_1164.all;		--�ޥήM��
Use IEEE.std_logic_unsigned.all;	--�ޥήM��

-- ----------------------------------------------------
entity Dht11_Driver is
	port(DHT11_CLK,DHT11_RESET:in std_logic;		--DHT11_CLK:781250Hz(50MHz/2^6:1.28us:FD(5))�ާ@�t�v,���m
		 DHT11_D_io:inout std_logic;				--DHT11 i/o
		 DHT11_DBo:out std_logic_vector(7 downto 0);--DHT11_driver ��ƿ�X
		 DHT11_RDp:in integer range 0 to 7;			--���Ū������
		 DHT11_tryN:in integer range 0 to 7;		--���~����մX��
		 DHT11_ok,DHT11_S:buffer std_logic;			--DHT11_driver�����@�~�X��,���~�H��
		 DHT11_DBoH,DHT11_DBoT:out integer range 0 to 255);--������X��פηū�
end entity Dht11_Driver;

-- -----------------------------------------------------
architecture Albert of Dht11_Driver is
	signal S_B,bit01,response:std_logic;	--start bit,�����줸
	signal ss:std_logic_vector(1 downto 0);	--���檬�A
	signal isdata:integer range 0 to 3;		--��ƪ��A
	signal dp,d8:integer range 0 to 7;		--��Ʀ줸�ާ@����
	signal dbit:std_logic_vector(6 downto 0);--byte
	signal chK_SUM:std_logic_vector(7 downto 0);--�d�M
	type DDataT is array(0 to 4) of std_logic_vector(7 downto 0);	--��ƽw�İϮ榡
	signal dd:DDataT;	--��ƽw�İ�
	signal tryNN:integer range 0 to 7;				--���~����մX��
	signal Timeout:std_logic_vector(21 downto 0);	--timeout�p�ɾ�
	signal tryDelay:integer range 0 to 31;
begin

DHT11_DBoH<=conv_integer(dd(4));--������X���(integer)
DHT11_DBoT<=conv_integer(dd(2));--������X�ū�(integer)

--DHT11_DBo��DHT11_RDp�����X��
DHT11_DBo<=dd(DHT11_RDp) when DHT11_RDp<5 else
		   chK_SUM 		 when DHT11_RDp=5 else (others=>'1');	--�W�Ǹ��

DHT11_D_io<='Z' when DHT11_RESET='0' or S_B='1' else '0';	--DHT11 data io �ާ@

DHT11:process(DHT11_CLK,DHT11_RESET)
begin
	if DHT11_RESET='0' then
		S_B<='0';				--start bit
		dp<=4;					--Ū��5byte
		d8<=7;					--Ū��8bit
		isdata<=2;				--��ƪ��A
		DHT11_ok<='0';			--�������@�~
		DHT11_S<='0';			--�Ѱ��@�~����
		tryNN<=DHT11_tryN;		--���~����մX��
		ss<="00";				--���檬�A��1�}�l
		Timeout<=(others=>'0');	--timeout�p�ɾ��k�s
		tryDelay<=11;			--11:��2.5ms,12:��5ms,13:��10ms,14:��21ms>18ms,15:��42ms>18ms
	elsif Rising_Edge(DHT11_CLK) and DHT11_ok='0' then
		Timeout<=Timeout+1;		--�p��
		case ss is
			----------------------------------------------------------
			--restart or Send request
			when "00"=>	--���� (restart:D_io->'Z')or(start bit:D_io->'0')
				if Timeout(tryDelay)='1' then	--start bit (�̦n��b2ms�H�W��í�w) Request DHT11
					tryDelay<=11;	--11:��2.5ms,12:��5ms,13:��10ms,14:��21ms,15:��42ms
					S_B<=not S_B;	--��X����줸
					Timeout<=(others=>'0');	--���_�p��
					ss<="0" & not S_B;		--���檬�A�U�@�B
					chK_SUM<=(others=>'0'); --�d�M�k�s
					response<='0';			--�U�ɤ��w���
				end if;

			----------------------------------------------------------
			--(Read response)
			--(Read each data segment and save it to a buffer)
			--end all stages

			--wait DHT11 Response pull low
			when "01"=>
				if DHT11_D_io='0' then
					Timeout<=(others=>'0');
					if isdata=0 then	--reciver bit
						d8<=d8-1;		--�������줸�ƻ���
						if d8=0 then	--�w����8bit
							dp<=dp-1;	--���������ƻ���
							dd(dp)<=dbit & bit01;	--�����줸�Φs�J��ƽw�İ�
							if dp<4 then
								chK_SUM<=chK_SUM+dd(dp+1); --�p��d�M
							end if;
							ss<="10";		--���檬�A�U�@�Bpull high
						else
							dbit<=dbit(5 downto 0) & bit01;--�����줸
							ss<="10";		--���檬�A�U�@�Bpull high
						end if;
					else
						isdata<=isdata-1;
						ss<="10";			--���檬�A�U�@�Bpull high
					end if;
				elsif Timeout=38 then		--��49us
					bit01<='1';				--�����줸0-->1
					--��Response(error)21ms>11~13ms	or DHT11 No data Response(error) --��164us
				elsif (Timeout(14)='1'and response='0')or(Timeout(7)='1'and response='1')  then
					ss<="11";				--���檬�A�U�@�B(���~�B�z)
				end if;		

			--wait DHT11 Response pull high
			when "10"=>
				if DHT11_D_io='1' then
					Timeout<=(others=>'0');	--���_�p��
					bit01<='0';				--�����줸�w�]0
					if dp=7 then --(�wŪ��40bit)stop bit
						if chK_SUM=dd(0) then
							DHT11_ok<='1';	--�@�~�w���T����
						else
							ss<="11";		--���檬�A�U�@�B(���~�B�z)
						end if;
					else
						ss<="01";			--���檬�A�U�@�B
					end if;
				elsif Timeout(7)='1' then	--DHT11 No Response(error) 7
					ss<="11";				--���檬�A�U�@�B(���~�B�z) --��164us
				end if;

			----------------------------------------------------------
			--"11"���~�B�z
			when others=>					--"11"���~�B�z
				if tryNN/=0 then
					tryNN<=tryNN-1;			--���տ��~�ƻ���
					Timeout<=(others=>'0');	--���_�p��
					dp<=4;					--����������
					d8<=7;					--�������줸��
					isdata<=2;				--�}�l���q
					tryDelay<=20;			--���Ȱ�1.4s
					ss<="00";				--restart
				else
					DHT11_ok<='1';			--�@�~�w����
					DHT11_S<='1';			--�@�~����
				end if;
		end case;
	end if;
end process;
--------------------------------------------
end Albert;