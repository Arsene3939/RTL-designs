--DM13A�X�ʾ�
--106.12.30��

Library IEEE;						--�s���s��w
Use IEEE.std_logic_1164.all;		--�ޥήM��
Use IEEE.std_logic_unsigned.all;	--�ޥήM��

-- ----------------------------------------------------
entity DM13A_Driver_RGB is
	port(--DM13A_Driver_RGB�ާ@�W�v,���m,ALE����,OE����,��V����,�Ϭ۱���
		 DM13ACLK,DM13A_RESET,DM13ALE,DM13AOE,BIT_R_L,not01:in std_logic;
		 startbit:in integer range 0 to 15;		 	--�}�l�ާ@�줸
		 maskRGB:in std_logic_vector(5 downto 0);	--�n�\�ާ@�줸
		 --mask (5):0:disable 1:enable, (4..3)00:load,01:xor:10:or,11:and RGB
		 LED_R,LED_G,LED_B:in std_logic_vector(15 downto 0);	--R G B �ϧΦ줸
		 DM13ACLKo,DM13ASDI_Ro,DM13ASDI_Go,DM13ASDI_Bo,DM13ALEo,DM13AOEo:out std_logic;--DM13A �w��ާ@�줸
		 DM13A_Sendok:out std_logic);	--DM13A_Driver_RGB�����ާ@�줸
end DM13A_Driver_RGB;

-- -----------------------------------------------------
architecture Albert of DM13A_Driver_RGB is
	signal DM13A_CLK:std_logic;					--DM13A CLK�����ާ@�줸
	signal i:integer range 0 to 31;				--��X�줸�Ʊ���
	constant databitN:integer range 0 to 31:=16;--��X�줸�ưѼ�:16 bit
	signal startbitS:integer range 0 to 15;		--�����}�l�ާ@�줸����
	signal R,G,B:std_logic;						--�����ϧΦ줸���X

-- --------------------------
begin

--R,G,B �ϧΦ줸���X�n�\�B��
R<=	LED_R(startbitS) when maskRGB(5)='0' else	--nop
	maskRGB(2)	 when BIT_R_L='1' and startbitS>startbit and maskRGB(4 downto 3)="00" else	--load
	maskRGB(2)	 when BIT_R_L='0' and startbitS<startbit and maskRGB(4 downto 3)="00" else	--load
	maskRGB(2) xor LED_R(startbitS)	 when BIT_R_L='1' and startbitS>startbit and maskRGB(4 downto 3)="01" else	--xor
	maskRGB(2) xor LED_R(startbitS)	 when BIT_R_L='0' and startbitS<startbit and maskRGB(4 downto 3)="01" else	--xor
	maskRGB(2) or  LED_R(startbitS)	 when BIT_R_L='1' and startbitS>startbit and maskRGB(4 downto 3)="10" else	--or
	maskRGB(2) or  LED_R(startbitS)	 when BIT_R_L='0' and startbitS<startbit and maskRGB(4 downto 3)="10" else	--or
	maskRGB(2) and LED_R(startbitS)	 when BIT_R_L='1' and startbitS>startbit and maskRGB(4 downto 3)="11" else	--and
	maskRGB(2) and LED_R(startbitS)	 when BIT_R_L='0' and startbitS<startbit and maskRGB(4 downto 3)="11" else	--and
	LED_R(startbitS);
G<=	LED_G(startbitS) when maskRGB(5)='0' else	--nop
	maskRGB(1)	 when BIT_R_L='1' and startbitS>startbit and maskRGB(4 downto 3)="00" else	--load
	maskRGB(1)	 when BIT_R_L='0' and startbitS<startbit and maskRGB(4 downto 3)="00" else	--load
	maskRGB(1) xor LED_G(startbitS)	 when BIT_R_L='1' and startbitS>startbit and maskRGB(4 downto 3)="01" else	--xor
	maskRGB(1) xor LED_G(startbitS)	 when BIT_R_L='0' and startbitS<startbit and maskRGB(4 downto 3)="01" else	--xor
	maskRGB(1) or  LED_G(startbitS)	 when BIT_R_L='1' and startbitS>startbit and maskRGB(4 downto 3)="10" else	--or
	maskRGB(1) or  LED_G(startbitS)	 when BIT_R_L='0' and startbitS<startbit and maskRGB(4 downto 3)="10" else	--or
	maskRGB(1) and LED_G(startbitS)	 when BIT_R_L='1' and startbitS>startbit and maskRGB(4 downto 3)="11" else	--and
	maskRGB(1) and LED_G(startbitS)	 when BIT_R_L='0' and startbitS<startbit and maskRGB(4 downto 3)="11" else	--and
	LED_G(startbitS);
B<=	LED_B(startbitS) when maskRGB(5)='0' else	--nop
	maskRGB(0)	 when BIT_R_L='1' and startbitS>startbit and maskRGB(4 downto 3)="00" else	--load
	maskRGB(0)	 when BIT_R_L='0' and startbitS<startbit and maskRGB(4 downto 3)="00" else	--load
	maskRGB(0) xor LED_B(startbitS)	 when BIT_R_L='1' and startbitS>startbit and maskRGB(4 downto 3)="01" else	--xor
	maskRGB(0) xor LED_B(startbitS)	 when BIT_R_L='0' and startbitS<startbit and maskRGB(4 downto 3)="01" else	--xor
	maskRGB(0) or  LED_B(startbitS)	 when BIT_R_L='1' and startbitS>startbit and maskRGB(4 downto 3)="10" else	--or
	maskRGB(0) or  LED_B(startbitS)	 when BIT_R_L='0' and startbitS<startbit and maskRGB(4 downto 3)="10" else	--or
	maskRGB(0) and LED_B(startbitS)	 when BIT_R_L='1' and startbitS>startbit and maskRGB(4 downto 3)="11" else	--and
	maskRGB(0) and LED_B(startbitS)	 when BIT_R_L='0' and startbitS<startbit and maskRGB(4 downto 3)="11" else	--and
	LED_B(startbitS);

--DM13A �w��ާ@�줸��X
DM13ASDI_Ro<=R xor not01;	--R SDI��X�B��(�Ϭ۱���)
DM13ASDI_Go<=G xor not01;	--G SDI��X�B��(�Ϭ۱���)
DM13ASDI_Bo<=B xor not01;	--B SDI��X�B��(�Ϭ۱���)
DM13ACLKo<=DM13A_CLK;		--CLK	
DM13ALEo<=DM13ALE;			--ALE
DM13AOEo<=DM13AOE;			--OE

DM13A_Send:process(DM13ACLK,DM13A_RESET)
begin
	if DM13A_RESET='0' then	--���m
		i<=0;				--��X�줸�ƭӼƹw�]0
		startbitS<=startbit;--���J�}�l�ާ@�줸
		DM13A_CLK<='0';		--�w�]Low
		DM13A_Sendok<='0';	--�w�]������
	elsif rising_edge(DM13ACLK) then
		if i=databitN then		--�P�_��X�줸�ƬO�_����
			DM13A_Sendok<='1';	--����
		else
			if DM13A_CLK='0' then
				DM13A_CLK<='1';	--�Ұʸ��JCLK
			else
				i<=i+1;			--��X�줸�Ƨ���1��
				DM13A_CLK<='0';	--�w�Ƹ��JCLK
				if BIT_R_L='1' then --���ˤ�V
					startbitS<=startbitS-1;	--�V�C�줸
				else
					startbitS<=startbitS+1;	--�V���줸
				end if;
			end if;
		end if;
	end if;
end process DM13A_Send;

--------------------------------------------
end Albert;
