--MCP4822 DAC����
--107.01.01��
--EP3C16Q240C8 50MHz LEs:15,408 PINs:161 ,gckp31 ,rstP99
--MCP4822_CH_BA:00(chA),01,11(chB),10->11(�۰ʥ�chA��chB:�����ഫ-�P�B��XDAC��) 

Library IEEE;						--�s���s��w
Use IEEE.std_logic_1164.all;		--�ޥήM��
Use IEEE.std_logic_unsigned.all;	--�ޥήM��
Use IEEE.std_logic_arith.all;		--�ޥήM��

-- ----------------------------------------------------
entity MCP4822_Driver is
	port(MCP4822_CLK,MCP4822_RESET:in std_logic;	--MCP4822_Driver�X��clk,reset�H��
		 MCP4822_DAA,MCP4822_DAB:in integer range 0 to 4095;	--MCP4822 DAC chA0,B1��
		 MCP4822_CHB_A:in std_logic_vector(1 downto 0);	--��J�q�D
		 MCP4822_GA_BA:in std_logic_vector(1 downto 0);	--GA 0x2,1x1
		 MCP4822_SHDN_BA:in std_logic_vector(1 downto 0);	--/SHDN
		 MCP4822_SDI,MCP4822_LDAC:out std_logic;		--MCP4822 SDI�H��
		 MCP4822_SCK,MCP4822_CS:buffer std_logic;		--MCP4822 SCK,/cs�H��
		 MCP4822_ok:buffer std_logic);	--Driver�����X�� ,�������A
end MCP4822_Driver;

-- -----------------------------------------------------
architecture Albert of MCP4822_Driver is
	signal i:integer range 0 to 15;			--�ާ@����
	signal MCP4822DAx,MCP4822DAB:std_logic_vector(14 downto 0);	--�ഫ��
	signal MCP4822_Chs:std_logic_vector(1 downto 0); 			--ch 0,1
-- --------------------------
begin

MCP4822:process(MCP4822_CLK,MCP4822_RESET)
begin
	if MCP4822_RESET='0' then		--���_�l:�ǳƸ��
		MCP4822_CS<='1';					--MCP4822 cs diable
		MCP4822_LDAC<='1';					--MCP4822 ldac diable
		MCP4822DAB<='0'&MCP4822_GA_BA(1)&MCP4822_SHDN_BA(1)&conv_std_logic_vector(MCP4822_DAB,12);		--B:DAC
		if MCP4822_CHB_A(0)='0' then
			MCP4822DAx<='0'&MCP4822_GA_BA(0)&MCP4822_SHDN_BA(0)&conv_std_logic_vector(MCP4822_DAA,12);	--A:DAC
		else
			MCP4822DAx<=MCP4822DAB;		--B:DAC
		end if;
		MCP4822_Chs<=MCP4822_CHB_A;			--�q�D���
		MCP4822_ok<='0';					--���m�ާ@�����X��
		i<=14;								--���m�ާ@����
	elsif rising_edge(MCP4822_CLK) then
		if MCP4822_ok='1' then				--�������ާ@
			MCP4822_LDAC<='1';					--����AC��
		elsif i=15 and MCP4822_SCK='1' then --write end
			MCP4822_CS<='1';					--MCP4822 cs diable
			MCP4822_Chs(0)<='1';				--chA-->chB�۰ʥ�chA��chB
			MCP4822DAx<=MCP4822DAB;				--B:DAC
			i<=14;								--�ǳƦ۰ʥ�chA��chB
			if MCP4822_Chs/="10" then			--����
				MCP4822_LDAC<='0';					--�ҰʷsAC��X
				MCP4822_ok<='1';					--�ާ@����
			end if;
		elsif MCP4822_CS='1' then			--���ާ@
			MCP4822_SDI<=MCP4822_Chs(0);		--CH bit
			MCP4822_CS<='0';					--enable /CS
			MCP4822_SCK<='0';					--���mMCP4822 /SCK
		else								--�ާ@��
			MCP4822_SCK<=not MCP4822_SCK;		--MCP4822 /SCK �ϦV
			if MCP4822_SCK='1' then	--clk H to L
				i<=i-1;							--�վ�ާ@����
				MCP4822_SDI<=MCP4822DAx(i);		--SDI out
			end if;
		end if;
	end if;
end process MCP4822;

--------------------------------------------
end Albert;
