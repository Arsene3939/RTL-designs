--Ws2812B RGB_LED�R�E�O2
--EP3C16Q240C8 50MHz LEs:15,408 PINs:161 ,gckP31 ,rstP99

Library IEEE;						--�s���s��w
Use IEEE.std_logic_1164.all;		--�ޥήM��
Use IEEE.std_logic_unsigned.all;	--�ޥήM��

entity CH3_WS2812B_2 is	
	port(gckP31,rstP99:in std_logic;--�t�έ��m�B�t�ήɯ�
		 WS2812Bout:out std_logic);	--WS2812B_Di�H����X(184)
end entity CH3_WS2812B_2;

architecture Albert of CH3_WS2812B_2 is
	--WS2812B�X�ʾ�------------------
	component WS2812B_Driver is
		port(	WS2812BCLK,WS2812BRESET,loadck:in std_logic;--�ާ@�W�v,���m,���Jck
				LEDGRBdata:in std_logic_vector(23 downto 0);--��m���
				reload,emitter,WS2812Bout:out std_logic		--�n�D���J,�o�g���A,�o�g��X 
			);
	end component;
	signal WS2812BCLK,WS2812BRESET,loadck,reload,emitter:std_logic;--�ާ@�W�v,���m,���Jck,�n�D���J,�o�g���A
	signal LEDGRBdata:std_logic_vector(23 downto 0);--��m���
	
	signal FD:std_logic_vector(24 downto 0);	--�t�ΰ��W��
	signal FD2:std_logic_vector(3 downto 0);	--WS2812B_Driver���W��
	signal SpeedS,WS2812BPCK:std_logic;			--WS2812BP�ާ@�W�v���,WS2812BP�ާ@�W�v
	signal delay:integer range 0 to 127;		--����ɶ�
	signal LED_WS2812B_N:integer range 0 to 127;--WS2812B�Ӽƫ���
	constant NLED:integer range 0 to 127:=29;	--WS2812B�Ӽ�:61��(0~60)
	signal LED_WS2812B_shiftN:integer range 0 to 7;--WS2812B����Ӽƫ���
	signal dir_LR:std_logic_vector(15 downto 0);   --��V����,WS2812BP�ާ@�W�v���,
	type LED_T is array(0 to 7) of std_logic_vector(23 downto 0);--�Ϲ��榡
	--�Ϲ�
	signal LED_WS2812B_T8:LED_T:=(--G       R       B
								"000000001111111100000000",
								"111111110000000000000000",
								"000000000000000011111111",
								"000000000000000000000000",
								"111111111111111100000000",
								"000000001111111111111111",
								"111111110000000011111111",
								"111111111111111111111111"
								);

begin

--WS2812B�X�ʾ�-----------------
WS2812BN: WS2812B_Driver port map(WS2812BCLK,WS2812BRESET,loadck,LEDGRBdata,reload,emitter,WS2812Bout);
		  WS2812BRESET<=rstP99;	--�t��reset

--��m��� ---------------------
LEDGRBdata<=LED_WS2812B_T8((LED_WS2812B_N+LED_WS2812B_shiftN) mod 8);

--WS2812BP�ާ@�W�v���
WS2812BPCK<=FD(8) when SpeedS='0' else 
			FD(16)when dir_LR(7)='0' else FD(18);--�̺C�t�v

WS2812BP:process(WS2812BPCK)
begin
	if rstP99='0' then
		LED_WS2812B_N<=0;	--�q�Y�}�l
		LED_WS2812B_shiftN<=0;--����0
		dir_LR<=(others=>'0');
		loadck<='0';
		SpeedS<='0';		--�[�־ާ@�t�v
	elsif rising_edge(WS2812BPCK) then
		if loadck='0' then	--���ݸ��J
			loadck<=reload;
		elsif LED_WS2812B_N=NLED then
			SpeedS<='1';			--��C�ާ@�t�v
			if emitter='0' then		--�w����o�g
				if delay/=0 then	--�I�G�ɶ�&�ܤƳt�v
					delay<=delay-1;	--�ɶ�����
				else
					loadck<='0';	--reemitter
					LED_WS2812B_N<=0;--�q�Y�}�l
					dir_LR<=dir_LR+1;--��V����
					if dir_LR(4)='1' then 
						LED_WS2812B_shiftN<=LED_WS2812B_shiftN+1;--���컼�W
					else
						LED_WS2812B_shiftN<=LED_WS2812B_shiftN-1;--���컼��
					end if;
					SpeedS<='0';	--�[�־ާ@�t�v
				end if;
			end if;
		else
			loadck<='0';
			LED_WS2812B_N<=LED_WS2812B_N+1;	--�վ��X��m
			delay<=20;
		end if;
	end if;
end process WS2812BP;

-- ���W��---------------------
Freq_Div:process(gckP31)
begin
	if rstP99='0' then		--�t�έ��m
		FD<=(others=>'0');
		FD2<=(others=>'0');
		WS2812BCLK<='0';			--WS2812BN�X���W�v
	elsif rising_edge(gckP31) then	--50MHz
		FD<=FD+1;					--���W��:2�i��W��(+1)�p�ƾ�
		if FD2=9 then				--7~12
			FD2<=(others=>'0');
			WS2812BCLK<=not WS2812BCLK;--50MHz/20=2.5MHz T.=. 0.4us
		else
			FD2<=FD2+1;				--���W��2:2�i��W��(+1)�p�ƾ�
		end if;
	end if;
end process Freq_Div;


end Albert;