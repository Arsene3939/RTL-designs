--LED�R�E�O1:�d��k
--EP3C16Q240C8 50MHz LEs:15,408 PINs:161 ,gckP31 ,rstP99

Library IEEE;						--�s���s��w
Use IEEE.std_logic_1164.all;		--�ޥήM��
Use IEEE.std_logic_unsigned.all;	--�ޥήM��

-- -----------------------------------------------------
entity CH2_LED_1 is
port(gckP31,rstP99:in std_logic;	-- �t�ήɯߡB�t�έ��m
	 LED16:buffer std_logic_vector(15 downto 0)	--LED
	 -- 87,93,95,94,100,101,102,103 
	 -- 106,107,108,110,111,112,113,114
	);
end entity CH2_LED_1; --or end CH2_LED_1;  --or end;

-- -----------------------------------------------------
architecture Albert of CH2_LED_1 is
	signal FD:std_logic_vector(24 downto 0);		--���W��
	type LED_T is array(0 to 127) of std_logic_vector(15 downto 0);--LED�˪O�榡
	constant LED_Tdata:LED_T:=	--LED�˪O���
	   (X"0000",X"8001",X"C003",X"E007",X"F00F",X"F81F",X"FC3F",X"FE7F",X"FFFF",X"7FFE",X"3FFC",X"1FF8",X"0FF0",X"07E0",X"03C0",X"0180",
		X"0000",X"0180",X"03C0",X"07E0",X"0FF0",X"1FF8",X"3FFC",X"7FFE",X"FFFF",X"FE7F",X"FC3F",X"F81F",X"F00F",X"E007",X"C003",X"8001",
		X"0000",X"0001",X"0005",X"0015",X"0055",X"0155",X"0555",X"1555",X"5555",X"5557",X"555F",X"557F",X"55FF",X"57FF",X"5FFF",X"7FFF",
		X"FFFF",X"BFFF",X"AFFF",X"ABFF",X"AAFF",X"AABF",X"AAAF",X"AAAB",X"AAAA",X"2AAA",X"0AAA",X"02AA",X"00AA",X"002A",X"000A",X"0002",
		X"0000",X"8001",X"C003",X"E007",X"F00F",X"F81F",X"FC3F",X"FE7F",X"FFFF",X"FE7F",X"FC3F",X"F81F",X"F00F",X"E007",X"C003",X"8001",
		X"0000",X"00FF",X"FF00",X"00FF",X"FF00",X"00FF",X"FF00",X"00FF",X"FF00",X"0000",X"FFFF",X"0000",X"FFFF",X"0000",X"FFFF",X"0000",
		X"FFFF",X"F00F",X"0FF0",X"F00F",X"0FF0",X"F00F",X"0FF0",X"F00F",X"0FF0",X"0000",X"0001",X"0003",X"0007",X"000F",X"001F",X"003F",
		X"007F",X"00FF",X"01FF",X"03FF",X"07FF",X"0FFF",X"1FFF",X"3FFF",X"7FFF",X"FFFF",X"0FFF",X"00FF",X"000F",X"0000",X"FFFF",X"0000");
	signal LED_T_p:integer range 0 to 127;		--LED_����
	signal LED_case:std_logic_vector(1 downto 0);	--����ﶵ

	signal PWM_reset:std_logic;--PWM�}��
	type PWM_T is array(0 to 15) of integer range 0 to 31;--PWM�榡
	signal LED_PWM:PWM_T;
	signal LED_PWM_data,not_LED:std_logic_vector(15 downto 0);--PWM,�Ϭ۱���

	signal speeds:integer range 0 to 3;	--�t�׿��
	signal speed:std_logic;				--����clk
	
-- --------------------------
begin

--LED��X�B��:	������				   �Ϭ�	  		 PWM
LED16<=(LED_Tdata(LED_T_p) xor not_LED) or LED_PWM_data;
--�t�׿ﶵ
speed<=FD(19) when speeds=0 else	--47.7Hz
	   FD(20) when speeds=1 else	--23.8Hz
	   FD(21) when speeds=2 else	--11.9Hz
	   FD(22);						--6Hz

--LED_P �D����----------------------------------------------
LED_P:process (speed,rstP99)
variable N:integer range 0 to 511;	--���榸��
variable LED_T_ps,LED_T_pe:integer range 0 to 127;	--�_�I,���I
variable dir_LR:std_logic;	--PWM��ʤ�V
begin
	if rstP99='0' then		--�t�έ��m
		N:=0;				--����ﶵ�w����
		LED_case<="00";		--����ﶵ�w�]
		speeds<=0;			--�t��0
	elsif rising_edge(speed) then
		if N=0 then	--����ﶵ�w����
			LED_case<=LED_case+1;	--����ﶵ�վ�
			case LED_case is		--����ﶵ�w�]��
				when "00"=>	
					N:=1;					--����ﶵ
					LED_T_p<=0;			--���Х�0�}�l
					LED_T_ps:=0;		--��0�}�l
					LED_T_pe:=127;	--��127����
					not_LED<=(others=>'0');	--���Ϭ�
					PWM_reset<='0';			--PWM off
				when "01"=>
					N:=1;					--����ﶵ
					LED_T_p<=0;			--���Х�0�}�l
					LED_T_ps:=0;		--��0�}�l
					LED_T_pe:=127;	--��127����
					not_LED<=(others=>'1');	--�Ϭ�
					PWM_reset<='0';			--PWM off
				when "10"=>
					N:=1;					--����ﶵ
					LED_T_p<=127;		--���Х�127�}�l
					LED_T_ps:=127;		--��127�}�l
					LED_T_pe:=0;		--��0����
					not_LED<=(others=>'0');	--���Ϭ�
					PWM_reset<='0';			--PWM off
				when "11"=>
					N:=127;					--����ﶵ
					LED_T_p<=0;			--���Х�0�}�l
					LED_T_ps:=0;		--��0�}�l
					LED_T_pe:=0;		--��0����
					not_LED<=(others=>'0');	--���Ϭ�
					dir_LR:='0';			--PWM��ʤ�V
					LED_PWM<=(0,0,1,2,3,4,5,7,10,12,15,17,20,24,28,31);
					--PWM�w�]��
					PWM_reset<='1';			--PWM on
					speeds<=speeds+1;		--�t�׽վ�
			end case;
		else	--����ﶵ
			if LED_T_ps=LED_T_pe then	--PWM�w�]�Ȳ���
				if dir_LR='0' then
					for i in 0 to 14 loop
						LED_PWM(i)<=LED_PWM(i+1);
					end loop;
					LED_PWM(15)<=LED_PWM(0);
				else
					for i in 0 to 14 loop
						LED_PWM(i+1)<=LED_PWM(i);
					end loop;
					LED_PWM(0)<=LED_PWM(15);
				end if;
				if (N mod 16)=0 then
					dir_LR:=not dir_LR;	--�վ�PWM��ʤ�V
				end if;
				N:=N-1;	--����-1
			elsif LED_T_ps<LED_T_pe then
				LED_T_p<=LED_T_p+1;	--���W
				if (LED_T_p+1)=LED_T_pe then
					N:=0;	--����
				end if;
			else
				LED_T_p<=LED_T_p-1;	--����
				if (LED_T_p-1)=LED_T_pe then
					N:=0;	--����
				end if;
			end if;
		end if;
	end if;
end process LED_P;

--PWM_P---------------------------------------------------
PWM_P:process(FD(0))
variable PWMc:integer range 0 to 31;	--PWM�p�ƾ�
begin
	if PWM_reset='0' then
		PWMc:=0;						--PWM�p�ƾ�
		LED_PWM_data<=(others=>'0');	--all on
	elsif rising_edge(FD(0)) then
		for i in 0 to 15 loop
			if LED_PWM(i)>PWMc then
				LED_PWM_data(i)<='0';	--on
			else
				LED_PWM_data(i)<='1';	--off
			end if;
		end loop;
		PWMc:= PWMc+1;					--PWM�p�ƾ��W��+1
	end if;
end process PWM_P;
	
-- ���W��----------------------------------------
Freq_Div:process(gckP31)			--�t���W�vgckP31:50MHz
begin
	if rstP99='0' then				--�t�έ��m
		FD<=(others=>'0');			--���W��:�k�s
	elsif rising_edge(gckP31) then	--50MHz
		FD<=FD+1;					--���W��:2�i��W��(+1)�p�ƾ�
	end if;
end process Freq_Div;

end Albert;
