--��I/O����
--EP3C16Q240C8 50MHz LEs:15,408 PINs:161 ,gckp31 ,SResetp99

library ieee;						--�s���s��w
use ieee.std_logic_1164.all;		--�ޥήM��
use ieee.std_logic_unsigned.all;	--�ޥήM��

entity ROTATE_ENCODER_EP3C16Q240C8 is 
--port(gckp31,SResetp99:in std_logic;				--�t���W�v,�t��reset
port(gckp31,ROTATEreset:in std_logic;				--�t���W�v,�t��reset
	 APi,BPi,PBi:in std_logic;
	 rsw:buffer std_logic_vector(2 downto 0)	--3�줸�p�ƾ�
	);
end ROTATE_ENCODER_EP3C16Q240C8;

architecture Albert of ROTATE_ENCODER_EP3C16Q240C8 is
	signal FD: std_logic_vector(25 downto 0);					--���W��
	signal APic,BPic,PBic:std_logic_vector(2 downto 0):="000";	--���u���p�ƾ�
begin

-- ����s�X�������q��----------------------------------------
EncoderInterface:process(APi,PBi,ROTATEreset)
begin
	if ROTATEreset='0' or PBic(2)='0' then	
		rsw<=(others=>'0');		-- �p�ƾ��k�s
	elsif rising_edge(APic(2)) then	-- ������UD�H�����ɽt��
		if BPi='1' then				-- �p�GB�H�������A�A�h�W��
			rsw<=rsw+1;
		else						-- �p�GB�H�����C�A�A�h�U��
			rsw<=rsw-1;
		end if;
	end if;
end process EncoderInterface; 

---------------------------------------------------------------
-- ���u���q��
Debounce:process(FD(8))	--����s�X�����u���W�v
begin

--APi���u���P���T
	if APi=APic(2) then	--�YAPi����APic�̥���줸
		APic<=APic(2) & "00";
		--�hAPi����APic(2)�k��줸�k�s
	elsif rising_edge(FD(8)) then	
		APic<=APic+1;
		--�_�h�HF1���ɽt�AAPic�p�ƾ����W
	end if;

--BPi���u���P���T
	if BPi=BPic(2) then	--�YBPi����BPic�̥���줸
		BPic<=BPic(2)& "00";	
		--�hBPi����BPic(2)�k��줸�k�s
	elsif rising_edge(FD(8)) then 
		BPic<=BPic+1;
		--�_�h�HF1���ɽt�ABPic�p�ƾ����W
	end if;

--PBi���u���P���T
	if PBi=PBic(2) then	--�YPBi����PBic�̥���줸
		PBic<=PBic(2)& "00";
		--�hPBic(2)�k��줸�k�s
	elsif rising_edge(FD(16)) then
		PBic<=PBic+1;
		--�_�h�HF1���ɽt�APBic�p�ƾ����W
	end if;
end process Debounce;

-- ���W��----------------------------------------
Freq_Div:process(GCKP31)
begin
	if ROTATEreset='0' then			--�t��reset
		FD<=(others=>'0');
	elsif rising_edge(GCKP31) then	--50MHz
		FD<=FD+1;
	end if;
end process Freq_Div;

end Albert;
