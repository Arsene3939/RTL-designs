--4��Ʊ��˦��@�����C�q��ܾ�
--�p�ƾ�:��ʭp�q��
--106.12.30��
--EP3C16Q240C8 50MHz LEs:15,408 PINs:161 ,gckp31 ,rstP99

Library IEEE;						--�s���s��w
Use IEEE.std_logic_1164.all;		--�ޥήM��
Use IEEE.std_logic_unsigned.all;	--�ޥήM��

-- ---------------------------------------
entity CH5_7SLED_1 is	
	port(gckP31,rstP99:in std_logic;--�t���W�v,�t��reset(�k�s)
		 S1,S8:in std_logic;		--���W���s(131),�k�s(117)
		 --4��Ʊ��y����ܾ�
		 SCANo:buffer std_logic_vector(3 downto 0);--���˾���X
		 Disp7S:buffer std_logic_vector(7 downto 0)--�p�Ʀ�ƸѽX��X
		 );
end entity CH5_7SLED_1;

-- -----------------------------------------
architecture Albert of CH5_7SLED_1 is
	signal FD:std_logic_vector(26 downto 0);	--�t�ΰ��W��
	type Disp7DataT is array(0 to 3) of integer range 0 to 9;--�p�ƾ��榡
	signal Disp7Data:Disp7DataT;				--�p�ƾ�
	signal scanP:integer range 0 to 3;			--���˾�����
	signal S1S,S8S:std_logic_vector(2 downto 0);--���u���p�ƾ�
begin

--�p�ƾ�--------------------------
counter_P:process(FD(18))
begin
	if rstP99='0' or S8S(2)='1' then	--�t�έ��m,�k�s
		Disp7Data(3)<=0;	--�p�ƾ�:�d���k�s
		Disp7Data(2)<=0;	--�p�ƾ�:�ʦ��k�s
		Disp7Data(1)<=0;	--�p�ƾ�:�Q���k�s
		Disp7Data(0)<=0;	--�p�ƾ�:�Ӧ��k�s
	elsif rising_edge(FD(18)) then
		if S1S(2)='1' then	--BCD�X���W
			if Disp7Data(0)/=9 then	Disp7Data(0)<=Disp7Data(0)+1; else Disp7Data(0)<=0;--�վ�Ӧ��
			if Disp7Data(1)/=9 then	Disp7Data(1)<=Disp7Data(1)+1; else Disp7Data(1)<=0;--�վ�Q���
			if Disp7Data(2)/=9 then	Disp7Data(2)<=Disp7Data(2)+1; else Disp7Data(2)<=0;--�վ�ʦ��
			if Disp7Data(3)/=9 then	Disp7Data(3)<=Disp7Data(3)+1; else Disp7Data(3)<=0;--�վ�d���
		end if;end if;end if;end if;end if;
	end if;
end process counter_P;

--4��Ʊ��˾�---------------------------------------------------
scan_P:process(FD(17),rstP99)
begin
	if rstP99='0' then
		scanP<=0;		--��ƨ��ȫ���
		SCANo<="1111";	--���˫H�� all off
	elsif rising_edge(FD(17)) then
		scanP<=scanP+1;	--��ƨ��ȫ��л��W
		SCANo<=SCANo(2 downto 0)&SCANo(3);
		if scanP=3 then		--�̫�@��ƤF
			scanP<=0;		----��ƨ��ȫ��Э��]
			SCANo<="1110";	--���˫H�����]
		end if;
	end if;
end process scan_P;

--BCD�X��:�@�����C�q��ܽXpgfedcba
with Disp7Data(scanP) select --���X��ܭ�
	Disp7S<=
	"11000000" when 0,
	"11111001" when 1,
	"10100100" when 2,
	"10110000" when 3,
	"10011001" when 4,
	"10010010" when 5,
	"10000010" when 6,
	"11111000" when 7,
	"10000000" when 8,
	"10010000" when 9,
	"11111111" when others;	--�����

----���u��----------------------------------
process(FD(17))
begin
	--S8���u��
	If S8='1' then
		S8S<="000";
	elsif rising_edge(FD(17)) then
		S8S<=S8S+ not S8S(2);
	end if;
	--S1���u��
	If S1='1' then
		S1S<="000";
	elsif rising_edge(FD(17)) then
		S1S<=S1S+ not S1S(2);
	end if;
end process;

-- --------------------------
--���W��
Freq_Div:process(gckP31)			--�t���W�vgckP31:50MHz
begin
	if rstP99='0' then				--�t�έ��m
		FD<=(others=>'0');			--���W��:�k�s
	elsif rising_edge(gckP31) then	--50MHz
		FD<=FD+1;					--���W��:2�i��W��(+1)�p�ƾ�
	end if;
end process Freq_Div;

-- ----------------------------------------
end Albert;