--LM35�ū׷P��������+MCP3202 ADC+����LCM���
--107.01.01��
--EP3C16Q240C8 50MHz LEs:15,408 PINs:161 ,gckp31 ,rstP99

Library IEEE;						--�s���s��w
Use IEEE.std_logic_1164.all;		--�ޥήM��
Use IEEE.std_logic_unsigned.all;	--�ޥήM��
Use IEEE.std_logic_arith.all;		--�ޥήM��

-- -----------------------------------------------------
entity CH11_LM35_ADC_1 is
port(gckP31,rstP99:in std_logic;--�t���W�v,�t��reset
	 --MCP3202
	 MCP3202_Di:out std_logic;
	 MCP3202_Do:in std_logic;
	 MCP3202_CLK,MCP3202_CS:buffer std_logic;
	 
	 --LCD 4bit����
	 DB_io:inout std_logic_vector(3 downto 0);
	 RSo,RWo,Eo:out std_logic
	 
	 );
end entity CH11_LM35_ADC_1;

-- -----------------------------------------------------
architecture Albert of CH11_LM35_ADC_1 is
	-- =ADC===========================================================================
	component MCP3202_Driver is
	port(MCP3202_CLK_D,MCP3202_RESET:in std_logic;	--MCP3202_Driver�X��clk,reset�H��
		 MCP3202_AD0,MCP3202_AD1:buffer integer range 0 to 4095;	--MCP3202 AD0,1 ch0,1��
		 MCP3202_try_N:in integer range 0 to 3;		--���ѫ�A���զ���
		 MCP3202_CH1_0:in std_logic_vector(1 downto 0);	--��J�q�D
		 MCP3202_SGL_DIFF:in std_logic;				--MCP3202 SGL/DIFF
		 MCP3202_Do:in std_logic;					--MCP3202 do�H��
		 MCP3202_Di:out std_logic;					--MCP3202 di�H��
		 MCP3202_CLK,MCP3202_CS:buffer std_logic;	--MCP3202 clk,/cs�H��
		 MCP3202_ok,MCP3202_S:buffer std_logic);	--Driver�����X�� ,�������A
	end component;
	
	signal MCP3202_CLK_D,MCP3202_RESET:std_logic;	--MCP3202_Driver�X��clk,reset�H��
	signal MCP3202_AD0,MCP3202_AD1:integer range 0 to 4095;--MCP3202 AD��
	signal MCP3202_try_N:integer range 0 to 3:=1;	--���ѫ�A���զ���
	signal MCP3202_CH1_0:std_logic_vector(1 downto 0):="01";--ch1
	signal MCP3202_SGL_DIFF:std_logic:='1';			--MCP3202 SGL/DIFF ��SGL
	signal MCP3202_ok,MCP3202_S:std_logic;			--Driver�����X�� ,�������A
			
	--------------------------------------------------------------------------------------
	--����LCM 4bit driver(WG14432B5)
	component LCM_4bit_driver is
	port(LCM_CLK,LCM_RESET:in std_logic;			--�ާ@�t�v,���m
		 RS,RW:in std_logic;						--�Ȧs�����,Ū�g�X�п�J
		 DBi:in std_logic_vector(7 downto 0);		--LCM_4bit_driver ��ƿ�J
		 DBo:out std_logic_vector(7 downto 0);		--LCM_4bit_driver ��ƿ�X
		 DB_io:inout std_logic_vector(3 downto 0);	--LCM DATA BUS����
		 RSo,RWo,Eo:out std_logic;					--LCM �Ȧs�����,Ū�g,�P�श��
		 LCMok,LCM_S:out boolean					--LCM_4bit_driver����,���~�X��
		 );
	end component;

	signal LCM_RESET,RS,RW:std_logic;				--LCM_4bit_driver���m,LCM�Ȧs�����,Ū�g�X��
	signal DBi,DBo:std_logic_vector(7 downto 0);	--LCM_4bit_driver�R�O�θ�ƿ�J�ο�X
	signal LCMok,LCM_S:boolean;						--LCM_4bit_driver�����@�~�X��,���~�H��

	-- ============================================================================
	signal FD:std_logic_vector(24 downto 0);--���W��
	signal times:integer range 0 to 2047;	--�p�ɾ�
	
	--------------------------------------------------------------
	----����LCM���O&��ƪ�榡:
	----(�`��,���O��,���O...���...........
	----�^�ƫ�LCM 4�줸�ɭ�,2�C���

	type LCM_T is array (0 to 20) of std_logic_vector(7 Downto 0);
	constant LCM_IT:LCM_T:=(X"0F",X"06",----���嫬LCM 4�줸�ɭ�
							"00101000","00101000","00101000",--4�줸�ɭ�
							"00000110","00001100","00000001",--ACC+1��ܹ��L����,��ܹ�on�L��еL�{�{,�M����ܹ�
							X"01",X"48",X"65",X"6C",X"6C",X"6F",X"21",X"20",X"20",X"20",x"20",X"20",X"20");--Hello!
	
	--LCM=1:�Ĥ@�C��ܰ�");-- -=MCP3202 ADC=-
	signal LCM_1:LCM_T:=(X"15",X"01",						--�`��,���O��
							"00000001",						--�M����ܹ�
							--��1�C��ܸ��
							X"20",X"2D",X"3D",X"4D",X"43",X"50",X"33",X"32",X"30",X"32",X"20",X"41",X"44",X"43",X"3D",X"2D",X"20",X"20");-- -=MCP3202 ADC=-

	--LCM=1:�ĤG�C��ܰ�LM35���ū׬�    �J
	signal LCM_12:LCM_T:=(X"15",X"01",						--�`��,���O��
							"10010000",						--�]�ĤG�CACC��m
							--��2�C��ܸ��
							X"4C",X"4D",X"33",X"35",X"B4",X"FA",X"B7",X"C5",X"AB",X"D7",X"AC",X"B0",X"20",X"20",X"20",X"20",X"A2",X"4A");--LM35���ū׬�    �J
	
	--LCM=2:�Ĥ@�C��ܰ�LM35 ���Ū������
	signal LCM_2:LCM_T:=(X"15",X"01",						--�`��,���O��
							"00000001",						--�M����ܹ�
							--��1�C��ܸ��
							X"4C",X"4D",X"33",X"35",X"20",X"20",X"B8",X"EA",X"AE",X"C6",X"C5",X"AA",X"A8",X"FA",X"A5",X"A2",X"B1",X"D1");--LM35 ���Ū������
	
	signal LCM_com_data,LCM_com_data2:LCM_T;--LCD����X
	signal LCM_INI:integer range 0 to 31;	--LCD����X����
	signal LCMP_RESET,LN,LCMPok:std_logic;	--LCM_P���m,��X�C��,LCM_P����
	signal LCM,LCMx:integer range 0 to 7;	--LCD��X�ﶵ
	
	signal lm35T:integer range 0 to 1550;	--LM35�ū׭�

-----------------------------
begin

U2: MCP3202_Driver port map(FD(4),MCP3202_RESET,		--MCP3202_Driver�X��clk,reset�H��
							MCP3202_AD0,MCP3202_AD1,	--MCP3202 AD��
							MCP3202_try_N,				--���ѫ�A���զ���
							MCP3202_CH1_0,				--��J�q�D
							MCP3202_SGL_DIFF,			--SGL/DIFF
							MCP3202_Do,					--MCP3202 do�H��
							MCP3202_Di,					--MCP3202 di�H��
							MCP3202_CLK,MCP3202_CS,		--MCP3202 clk,/cs�H�� 
							MCP3202_ok,MCP3202_S);		--Driver�����X�� ,�������A
--����LCM				  
LCMset: LCM_4bit_driver port map(FD(7),LCM_RESET,RS,RW,DBi,DBo,DB_io,RSo,RWo,Eo,LCMok,LCM_S);	--LCM�Ҳ�

-----------------------------
LM35P_Main:process(FD(17))
begin
	if rstP99='0' then			--�t�έ��m
		MCP3202_RESET<='0';		--MCP3202_Driver off
		LCM<=0;					--����LCM��l��
		LCMP_RESET<='0';		--LCMP���m
	elsif rising_edge(FD(17)) then
		LCMP_RESET<='1';		--LCMP�Ұ����	
		if LCMPok='1' then
			if MCP3202_RESET='0' then	--MCP3202_Driver�|���Ұ�
				MCP3202_RESET<='1';		--ADC���Ū��
				times<=400;				--�]�w�p��
			elsif MCP3202_ok='1' then	--ADCŪ������
				times<=times-1;			--�p��
				if times=0 then			--�ɶ���
					LCM<=1;				--����LCM��ܴ��q��
					LCMP_RESET<='0';	--LCMP���m
					MCP3202_RESET<='0';	--MCP3202_Driver�ǳƭ��sŪ�����
				elsif MCP3202_S='1' then--���Ū������
					LCM<=2;				--����LCM��� LM35 ���Ū������
				end if;
			end if;
		end if;
	end if;
end process LM35P_Main;

------------------------------------------------------------
--LM35:LCM���
LM35T<=MCP3202_AD1*122/100;	--5/10mv=500/4095*1000=122*MCP3202_AD1/100
LCM_12(18)<="0011" & conv_std_logic_vector(LM35T mod 10,4);			-- �^���p��1��
LCM_12(17)<=X"2E";													--.�p���I
LCM_12(16)<="0011" & conv_std_logic_vector((LM35T/10) mod 10,4);	-- �^���Ӧ��
LCM_12(15)<="0011" & conv_std_logic_vector(LM35T/100,4);			-- �^���Q���

--�[��ADC�ഫ��X
--LCM_12(18)<="0011" & conv_std_logic_vector(MCP3202_AD1 mod 10,4);		-- �^���Ӧ��
--LCM_12(17)<="0011" & conv_std_logic_vector((MCP3202_AD1/10)mod 10,4);	-- �^���Q���
--LCM_12(16)<="0011" & conv_std_logic_vector((MCP3202_AD1/100) mod 10,4);	-- �^���ʦ��
--LCM_12(15)<="0011" & conv_std_logic_vector(MCP3202_AD1/1000,4);			-- �^���d���

--����LCM��ܾ�---------------------------------------------------
--����LCM��ܾ�
--���O&��ƪ�榡: 
--(�`��,���O��,���O...���..........
LCM_P:process(FD(0))
	variable SW:Boolean;				--�R�O�θ�ƳƧ��X��
begin
	if LCM/=LCMx or LCMP_RESET='0' then
		LCMx<=LCM;						--�O���ﶵ
		LCM_RESET<='0';					--LCM���m
		LCM_INI<=2;						--�R�O�θ�Ư��޳]���_�I
		LN<='0';						--�]�w��X1�C
		case LCM is
			when 0=>
				LCM_com_data<=LCM_IT;	--LCM��l�ƿ�X�Ĥ@�C���Hello!
			when 1=>
				LCM_com_data<=LCM_1;	--��X�Ĥ@�C���
				LCM_com_data2<=LCM_12;	--��X�ĤG�C���
				LN<='1';				--�]�w��X2�C
			when others =>
				LCM_com_data<=LCM_2;	--��X�Ĥ@�C���
		end case;
		LCMPok<='0';					--���������H��
		SW:=False;						--�R�O�θ�ƳƧ��X��
	elsif rising_edge(FD(0)) then
		if SW then						--�R�O�θ�ƳƧ���
			LCM_RESET<='1';				--�Ұ�LCM_4bit_driver_delay
			SW:=False;					--���m�X��
		elsif LCM_RESET='1' then		--LCM_4bit_driver_delay�Ұʤ�
			if LCMok then				--����LCM_4bit_driver_delay�����ǰe
				LCM_RESET<='0';			--������LCM���m
			end if;
		elsif LCM_INI<LCM_com_data(0) and LCM_INI<LCM_com_data'length then	--�R�O�θ�Ʃ|���ǧ�
			if LCM_INI<=(LCM_com_data(1)+1) then--��R�O�θ�ƼȦs��
				RS<='0';	--Instruction reg
			else
				RS<='1';	--Data reg
			end if;
			RW<='0';		--LCM�g�J�ާ@
			DBi<=LCM_com_data(LCM_INI);	--���J�R�O�θ��
			LCM_INI<=LCM_INI+1;			--�R�O�θ�Ư��ޫ���U�@��
			SW:=True;					--�R�O�θ�Ƥw�Ƨ�
		else
			if LN='1' then				--�]�w��X2�C
				LN<='0';					--�]�w��X2�C����
				LCM_INI<=2;					--�R�O�θ�Ư��޳]���_�I
				LCM_com_data<=LCM_com_data2;--LCM��X�ĤG�C���
			else
				LCMPok<='1';				--���槹��
			end if;
		end if;
	end if;
end process LCM_P;	

----���W��--------------------------
Freq_Div:process(gckP31)			--�t���W�vgckP31:50MHz
begin
	if rstP99='0' then				--�t�έ��m
		FD<=(others=>'0');			--���W��:�k�s
	elsif rising_edge(gckP31) then	--50MHz
		FD<=FD+1;					--���W��:2�i��W��(+1)�p�ƾ�
	end if;
end process Freq_Div;

-- ----------------------------------------
end Albert;
