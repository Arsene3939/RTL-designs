--MCP3202 ADC����
--107.01.01��
--EP3C16Q240C8 50MHz LEs:15,408 PINs:161 ,gckp31 ,rstP99
--MCP3202: MSBF='1'
--MCP3202_CH1_0:00(ch0),01,11(ch1),10->11(�۰ʥ�ch0��ch1:�����ഫ-�P�B��XADC��) 

Library IEEE;						--�s���s��w
Use IEEE.std_logic_1164.all;		--�ޥήM��
Use IEEE.std_logic_unsigned.all;	--�ޥήM��

-- ----------------------------------------------------
entity MCP3202_Driver is
	port(MCP3202_CLK_D,MCP3202_RESET:in std_logic;	--MCP3202_Driver�X��clk,reset�H��
		 MCP3202_AD0,MCP3202_AD1:buffer integer range 0 to 4095;	--MCP3202 AD0,1 ch0,1��
		 MCP3202_try_N:in integer range 0 to 3;		--���ѫ�A���զ���
		 MCP3202_CH1_0:in std_logic_vector(1 downto 0);	--��J�q�D
		 MCP3202_SGL_DIFF:in std_logic;				--MCP3202 SGL/DIFF
		 MCP3202_Do:in std_logic;					--MCP3202 do�H��
		 MCP3202_Di:out std_logic;					--MCP3202 di�H��
		 MCP3202_CLK,MCP3202_CS:buffer std_logic;	--MCP3202 clk,/cs�H��
		 MCP3202_ok,MCP3202_S:buffer std_logic);	--Driver�����X�� ,�������A
end entity MCP3202_Driver;

-- -----------------------------------------------------
architecture Albert of MCP3202_Driver is
	signal MCP3202_tryN:integer range 0 to 3;		--���ѫ�A���զ���
	signal MCP3202Dis:std_logic_vector(2 downto 0);	--2:MSBF+1:ODD/SIGN+0:SGL/DIFF
	signal MCP3202_ADs:std_logic_vector(11 downto 0);--�ഫ�Ȧ���
	signal MCP3202_Chs:std_logic_vector(1 downto 0); --ch 0,1
	signal i:integer range 0 to 31;					--�ާ@����
-- --------------------------
begin

MCP3202:process(MCP3202_CLK_D,MCP3202_RESET)
begin
	if MCP3202_RESET='0' then		--���_�l
		MCP3202_CS<='1';					--MCP3202 cs diable
		MCP3202_tryN<=MCP3202_try_N;		--���ѫ�A���զ���(�_�l��L�k�A��)
		MCP3202_Chs<=MCP3202_CH1_0;			--�q�D���(�_�l��L�k�A��)
		MCP3202_ok<='0';					--���m�ާ@�����X��
		MCP3202_S<='0';						--���m�������A
		MCP3202Dis<='1'&MCP3202_CH1_0(0)&MCP3202_SGL_DIFF;	--2:MSBF+1:ODD/SIGN+0:SGL/DIFF(�_�l��L�k�A��)
	elsif rising_edge(MCP3202_CLK_D) then
		if MCP3202_ok='0' then		--�������ާ@
			if i=17 then 				--read end
				if MCP3202Dis(1)='0' then
					MCP3202_AD0<=conv_integer(MCP3202_ADs);	--ch0 ADC��
				else
					MCP3202_AD1<=conv_integer(MCP3202_ADs);	--ch1 ADC��
				end if;
				i<=0;						--���m�ާ@����
				MCP3202_CS<='1';			--MCP3202 cs diable
				MCP3202Dis(1)<='1';			--ch0-->ch1
				MCP3202_ok<=not MCP3202_Chs(1) or MCP3202Dis(1);--�۰ʥ�ch0��ch1 or �ާ@����,���\����
			elsif MCP3202_CS='1' then	--���ާ@
				i<=0;						--���m�ާ@����
				MCP3202_Di<='1';				--start bit
				MCP3202_CS<='0';			--enable /CS
				MCP3202_CLK<='0';			--���mMCP3202 /CLK
			else						--�ާ@��
				MCP3202_CLK<=not MCP3202_CLK;--MCP3202 /CLK �ϦV
				if MCP3202_CLK='1' then	--clk H to L:Di out
					if i<3 then				--MCP3202 �_�l���q
						MCP3202_Di<=MCP3202Dis(i);	--2:MSBF+1:ODD/SIGN+0:SGL/DIFF
						i<=i+1;				--�վ�ާ@����
					end if;
				elsif i>2 then			--clk L to H:Do in --�i�J�������q
					i<=i+1;					--�վ�ާ@����
					MCP3202_ADs<=MCP3202_ADs(10 downto 0)&MCP3202_Do;--�ഫ�Ȧ���
					if i=4 and MCP3202_Do='1' then --error
						MCP3202_tryN<=MCP3202_tryN-1;	--���ѫ�վ�A���զ���
						if MCP3202_tryN=0 then	--���Ѥ��ΦA�դF
							MCP3202_ok<='1';	--�ާ@����
							MCP3202_S<='1';		--����
						else			--retry
							MCP3202_CS<='1';--MCP3202 cs diable
						end if;
					end if;
				end if;
			end if;
		end if;
	end if;
end process MCP3202;

--------------------------------------------
end Albert;
