--DoReMi�B����IC ����
--107.01.01��
--EP3C16Q240C8 50MHz LEs:15,408 PINs:161 ,gckp31 ,rstP99

Library IEEE;						--�s���s��w
Use IEEE.std_logic_1164.all;		--�ޥήM��
Use IEEE.std_logic_unsigned.all;	--�ޥήM��

-- ----------------------------------------------------
entity CH8_SOUND_1 is
	Port(gckP31,rstP99:in std_logic;--�t���W�v,�t��reset
		 S1,S2:in std_logic;		--����IC���s�B�~�E�����ﾹ���s
		 --����IC�B�~�E�����ﾹ��X
		 MusicIC,Do_Re_Mio:out std_logic
		 );
end entity CH8_SOUND_1;

-- ----------------------------------------------------
architecture Albert of CH8_SOUND_1 is
	--DoReMi_S Driver----------------------------------
	component DoReMi_S is
	Port(CLK,Sound_RESET,S_P_N:in std_logic;	--�t�ήɯ�,�t�έ��m
		 ToneS:in integer range 0 to 37;		--����
		 BeatS:in std_logic_vector(9 downto 0);	--�`��
		 Soundend,Do_Re_Mio:out std_logic);		--������,����X
	end component;

	signal Sound_RESET,Soundend:std_logic;--���m,������
	signal S_WAIT:integer range 0 to 3;			 --���ݭ�����
	signal BeatS:std_logic_vector(9 downto 0);	 --�`��
	signal ToneS:integer range 0 to 37;			 --����

	---------------------------------------------------
	signal FD:std_logic_vector(24 downto 0);	--���W��
	signal UpDn,S_L_UD:std_logic;				--�ɭ������B�`��
	signal S_L:std_logic_vector(4 downto 0);	--�`��վ㭿�v
	signal S1S,S2S:std_logic_vector(2 downto 0);--���u���p�ƾ�
	signal MusicIC_on,Sound_main_reset,S2_off:std_logic:='0';--����IC��X����,Sound_main���m,S2����
	
begin

--DoReMi_S Driver--------------------------------------------
U1: DoReMi_S port map(gckp31,Sound_RESET,'1',ToneS,BeatS,Soundend,Do_Re_Mio);

MusicIC<=MusicIC_on;--S1S(2);--����IC��X

--�`��--------------------------------------------
BeatS<="0000001010" + S_L * "00101";	--0.1s~1.65s�`��վ�

--���s�ާ@------------------------------------
process(FD(18))
begin
	--����IC���s
	if rising_edge(FD(18)) then
		if S1S(2)='1' then
			--����IC��X����
			MusicIC_on<=not MusicIC_on;
		end if;
	end if;
	--�~�E�����ﾹ���s
	if S2S=0 then					--S2���s��}
		Sound_main_reset<=S2_off;	--Sound_main on_off����
	elsif rising_edge(FD(18)) then
		if S2S(2)='1' then
			--Sound_main on_off����
			Sound_main_reset<=not Sound_main_reset;
		end if;
	end if;
end process;

--Sound_main-----------------------------------------
Sound_main:process(FD(0))
begin
	if Sound_main_reset='0' then
		ToneS<=0;			--�����w�]:0
		S_L<="00000";		--�`��վ㭿�v�w�]:0
		UpDn<='1';			--�ɭ������w�]:��
		S_L_UD<='1';		--�ɭ��`��w�]:��
		Sound_RESET<='0';	--DoReMi_S���m
		S2_off<='0';		--����Sound_main_reset
	elsif rising_edge(FD(0)) then
		if S_L/="10000" then
			S2_off<='1';			--�����Ұ�Sound_main_reset
			if Soundend='1' then	--DoReMi_S �������F
				Sound_RESET<='0';	--DoReMi_S���m
				if UpDn='1' then	--�ɭ���
					ToneS<=ToneS+1;	--�ɭ���
					if ToneS=36 then--�̰��@�ӤF
						UpDn<='0';	--�ﭰ����
					end if;
				else	--������
					ToneS<=ToneS-1;			--������
					if ToneS=1 then			--�̧C�@�ӤF
						UpDn<='1';			--��ɭ���
						if S_L_UD='1' then	--�ɸ`��(�[��)
							S_L<=S_L+1;		--�[��
							if S_L=3 then	--�̪��F
								S_L_UD<='0';--�ﭰ�`��(�ܵu)
							end if;
						else				--���`��
							S_L<=S_L-1;		--�ܵu
							if S_L=1 then	--�̵u�F
								--Sound_main�����F
								S_L<="10000";--��S2���s����}
								--�^��Sound_main_reset
								S2_off<='0';
							end if;
						end if;
					end if;
				end if;
			else
				Sound_RESET<='1';	--�Ұ�DoReMi_S
			end if;
		end if;
	end if;
end process Sound_main;

--���u��----------------------------------
process(FD(17))
begin
	--S1���u��--����IC���s
	if S1='1' then
		S1S<="000";
	elsif rising_edge(FD(17)) then
		S1S<=S1S+ not S1S(2);
	end if;
	--S2���u��--�~�E�����ﾹ���s
	if S2='1' then
		S2S<="000";
	elsif rising_edge(FD(17)) then
		S2S<=S2S+ not S2S(2);
	end if;
end process;

----���W��--------------------------
Freq_Div:process(gckP31)			--�t���W�vgckP31:50MHz
begin
	if rstP99='0' then				--�t�έ��m
		FD<=(others=>'0');			--���W��:�k�s
	elsif rising_edge(gckP31) then	--50MHz
		FD<=FD+1;					--���W��:2�i��W��(+1)�p�ƾ�
	end if;
end process Freq_Div;

-- ----------------------------------------
end Albert;