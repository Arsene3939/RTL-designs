--DHT11����׷P��������:1 wire
--107.01.01��
--EP3C16Q240C8 50MHz LEs:15,408 PINs:161 ,gckp31 ,rstP99

Library IEEE;						--�s���s��w
Use IEEE.std_logic_1164.all;		--�ޥήM��
Use IEEE.std_logic_unsigned.all;	--�ޥήM��
Use IEEE.numeric_std.all;			--�ޥήM��

-- -----------------------------------------------------
entity CH10_DHT11_2 is
port(gckP31,rstP99:in std_logic;--�t���W�v,�t��reset
     sw8_1,sw8_2:in std_logic_vector(7 downto 0);	--�����}����J:�ū׳]�w,��׳]�w
	 --DHT11
	 DHT11_D_io:inout std_logic;	--DHT11 i/o
	 
	 --DHT11 �C�q��ܾ���ܿ�X
	 DHT11_scan:buffer unsigned(3 downto 0);	--���˫H��
	 D7data:out std_logic_vector(7 downto 0);	--��ܸ��
	 D7xx_xx:out std_logic;	--:
	 
	 --���ﾹ��X
	 sound1,sound2:buffer std_logic
    );
end entity CH10_DHT11_2;

-- -----------------------------------------------------
architecture Albert of CH10_DHT11_2 is
	-- ============================================================================
	--DHT11_driver
	--Data format:
	--DHT11_DBo(std_logic_vector:8bit):��DHT11_RDp�����X��
	--RDp=5:chK_SUM
	--RDp=4							   3							   2								1								  0					
	--The 8bit humidity integer data + 8bit the Humidity decimal data +8 bit temperature integer data + 8bit fractional temperature data +8 bit parity bit.
	--������X���(DHT11_DBoH)�ηū�(DHT11_DBoT):integer(0~255:8bit)
	--105.11.30��
	component DHT11_driver is
		port(DHT11_CLK,DHT11_RESET:in std_logic;		--DHT11_CLK:781250Hz(50MHz/2^6:1.28us:FD(5))�ާ@�t�v,���m
			 DHT11_D_io:inout std_logic;				--DHT11 i/o
			 DHT11_DBo:out std_logic_vector(7 downto 0);--DHT11_driver ��ƿ�X
			 DHT11_RDp:in integer range 0 to 7;			--���Ū������
			 DHT11_tryN:in integer range 0 to 7;		--���~����մX��
			 DHT11_ok,DHT11_S:buffer std_logic;			--DHT11_driver�����@�~�X��,���~�H��
			 DHT11_DBoH,DHT11_DBoT:out integer range 0 to 255);--������X��פηū�
	end component DHT11_driver;
	signal DHT11_CLK,DHT11_RESET:std_logic;	--DHT11_CLK:781250Hz(50MHz/2^6:1.28us:FD(5))�ާ@�t�v,���m
	signal DHT11_DBo:std_logic_vector(7 downto 0);--DHT11_driver ��ƿ�X
	signal DHT11_RDp:integer range 0 to 7;		--���Ū������5~0
	signal DHT11_tryN:integer range 0 to 7:=3;	--���~����մX��
	signal DHT11_ok,DHT11_S:std_logic;			--DHT11_driver�����@�~�X��,���~�H��	
	signal DHT11_DBoH,DHT11_DBoT:integer range 0 to 255;--������X��פηū�

	-- ============================================================================
	signal FD:std_logic_vector(24 downto 0);--���W��
	signal scanP:integer range 0 to 3;		--��ƨ��ȫ���
	signal HL,TL:std_logic;					--��סB�ūת��A
	signal D7sp:std_logic;					--�p���I
	signal Disp7S:std_logic_vector(6 downto 0);	--��ܸѽX

	type D7_data_T is array (0 to 3) of integer range 0 to 15;--DHT11��ܭȮ榡
	signal D7_data:D7_data_T:=(0,0,0,0);	--DHT11��ܭ�
	signal times:integer range 0 to 2047;	--�p�ɾ�

begin
-----------------------------
DHT11_CLK<=FD(5);	--DHT11_CLK:781250Hz(50MHz/2^6:1.28us:FD(5))�ާ@�t�v
U2: DHT11_driver port map(DHT11_CLK,DHT11_RESET,--DHT11_CLK:781250Hz(50MHz/2^6:1.28us:FD(5))�ާ@�t�v,���m
						  DHT11_D_io,			--DHT11 i/o
						  DHT11_DBo,			--DHT11_driver ��ƿ�X
						  DHT11_RDp,			--���Ū������
						  DHT11_tryN,			--���~����մX��
						  DHT11_ok,DHT11_S,DHT11_DBoH,DHT11_DBoT);	--DHT11_driver�����@�~�X��,���~�H��,������X��פηū�

-----------------------------
DHT11P_Main:process(FD(17))
begin
	if rstP99='0' then	--�t�έ��m
		DHT11_RESET<='0';		--DHT11�ǳƭ��sŪ�����
		D7xx_xx<='1';			--:���G
	elsif rising_edge(FD(17)) then
		if DHT11_RESET='0' then	--DHT11_driver�|���Ұ�
			DHT11_RESET<='1';		--DHT11���Ū��
			D7xx_xx<='0';			--:�G (DHT11���Ū��)
			times<=1400;			--�]�w�p��
		elsif DHT11_ok='1' then	--DHT11Ū������
			D7xx_xx<='1';			--:���G (DHT11Ū������)
			times<=times-1;			--�p��
			if times=0 then		--�ɶ���
				DHT11_RESET<='0';	--DHT11�ǳƭ��sŪ�����
			end if;
		end if;
	end if;
end process DHT11P_Main;

------------------------------------------------------------
--���ﾹ��X
--���ĵ���n
HL<='0' when DHT11_DBoH>(conv_integer(sw8_2(7 downto 4))*10+conv_integer(sw8_2(3 downto 0))) else '1';
sound1<=FD(22)and FD(16)and not HL;
--�ū�ĵ���n
TL<='0' when DHT11_DBoT>(conv_integer(sw8_1(7 downto 4))*10+conv_integer(sw8_1(3 downto 0))) else '1';
sound2<=not TL;

--DHT11 ���
D7_data(0)<=DHT11_DBoH mod 10;		-- ����^���Ӧ��
D7_data(1)<=(DHT11_DBoH/10)mod 10;	-- ����^���Q���
D7_data(2)<=DHT11_DBoT mod 10;		-- �ū��^���Ӧ��
D7_data(3)<=(DHT11_DBoT/10)mod 10;	-- �ū��^���Q���

--4��Ʊ��˾�----------------------------------------
scan_P:process(FD(17))
begin
	if rstP99='0' then
		scanP<=0;		--��ƨ��ȫ���
		DHT11_scan<="1111";	--���˫H��
	elsif rising_edge(FD(17)) then
		scanP<=scanP+1;
		DHT11_scan<=DHT11_scan rol 1; --DHT11_scan ������unsigned
		--DHT11_scan<=DHT11_scan(2 downto 0) & DHT11_scan(3);-- DHT11_scan �i��unsigned��std_logic_vector
		if scanP=3 then
			scanP<=0;
			DHT11_scan<="1110";	--���˫H��
		end if;
	end if;
end process scan_P;

--�p���I����(�{�{��ܶW�X�]�w)
with scanP select
	D7sp<=
	HL when 0,--���
	HL when 1,--���
	TL when 2,--�ū�
	TL when 3;--�ū�

D7data<=(D7sp or FD(24)) & Disp7S;--�C�q��ܽX��X��X

--BCD�X�Ѧ@�����C�q��ܽXpgfedcba
with D7_data(scanP) select --���X��ܭ�
	Disp7S<=
	"1000000" when 0,
	"1111001" when 1,
	"0100100" when 2,
	"0110000" when 3,
	"0011001" when 4,
	"0010010" when 5,
	"0000010" when 6,
	"1111000" when 7,
	"0000000" when 8,
	"0010000" when 9,
	"1111111" when others;	--�����

----���W��--------------------------
Freq_Div:process(gckP31)			--�t���W�vgckP31:50MHz
begin
	if rstP99='0' then				--�t�έ��m
		FD<=(others=>'0');			--���W��:�k�s
	elsif rising_edge(gckP31) then	--50MHz
		FD<=FD+1;					--���W��:2�i��W��(+1)�p�ƾ�
	end if;
end process Freq_Div;

-- ----------------------------------------
end Albert;
