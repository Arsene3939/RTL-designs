--2017.04.30��(V2)
--EP3C16Q240C8 50MHz LEs:15,408 PINs:161 ,gckp31 ,SResetp99
--Bluetooth_UART ����+PC+����LCM���
--BT_RX=147, BT_TX=148
--USB_RX=144,USB_TX=145

--on=0�Boff=1
--DIP1 
-- on(0)  ������
-- off(1) �۰ʤ���0~7
--DIP2�BDIP3
-- on(0)�Bon(0)	�G��DIP6,DIP7,DIP8��������
-- on(0)�Boff(1)�G�� ����s�X�� ��������
-- off(1)�Bon(0)�G�� ��L0~7 ��������
-- off(1)�Boff(1)�G�� �Ť�/USB ��������

--DIP6�BDIP7�BDIP8:
--0:000:����
--1:001:LED16�q
--2:010:���ﾹ��X
--3:011:DHT11 ����״��� (�W�� DHT11 ��,���:2byte)
--4:100:WS2812B test
--5:101:MG90S test.
--6:110:RGB16x16 test
--7:111:LM35 test (�W�� ADC:2byte)
--����:S7�ծ�S8�դ�

--dip15P57�G����USB/BT
--on(0)USB�Boff(1)BT 

--dip16P56�G�s�򼽩�ɤ��n���}��
--on(0)����Boff(1)�R�� 

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

-- -----------------------------------------------------
entity KTM626 is
port(GCKP31,SResetP99:in std_logic;		--�t���W�v,�t��reset
	s0,s1,s2,M0,M1,M2:in std_logic;		--�ާ@�����}��
	--UART BT
--	BT_RX:in std_logic;		--RD=BT_RX
--	BT_TX:out std_logic;	--TX=BT_TX
	--UART USB
--	USB_RX:in std_logic;
--	USB_TX:out std_logic;

	--UART BT(����)
	BT_RX:out std_logic;
	BT_TX:in std_logic;	
	--UART USB(����)
	USB_RX:out std_logic;
	USB_TX:in std_logic;

	dip15P57:in std_logic;	--on(0)=USB, off(1)=BT
	
	--DHT11 i/o
	DHT11_D_io:inout std_logic;
	--LCD 4bit����
	DB_io:inout std_logic_vector(3 downto 0);
	RSo,RWo,Eo:out std_logic;
	--LED16�q
	led16:buffer std_logic_vector(15 downto 0);
	--���ﾹ��X
	sound1,sound2:buffer std_logic;
	dip16P56:in std_logic;
	--��C��LED�H����X
	WS2812Bout:out std_logic;
	--MG90S���A����X
	MG90S_o0:out std_logic;
	MG90S_o1:out std_logic;
	--RGB16x16��X
	DM13ACLKo,DM13ASDI_Ro,DM13ASDI_Go,DM13ASDI_Bo,DM13ALEo,DM13AOEo:out std_logic;
	Scan_DCBAo:buffer std_logic_vector(3 downto 0);
	--MCP3202 ADC
	MCP3202_Di:out std_logic;
	MCP3202_Do:in std_logic;
	MCP3202_CLK,MCP3202_CS:buffer std_logic;
	--timer0�Ʀ����
	PB7,PB8: in std_logic;					--�ծ�,�դ����s
	scan:buffer unsigned(3 downto 0);			--���˫H��
	D7data:out std_logic_vector(6 downto 0);	--��ܸ��
	D7xx_xx:out std_logic;					--:�{��
	--����s�X��_���
	APi,BPi,PBi:in std_logic;
	--��L_���
	keyi:in std_logic_vector(3 downto 0);		--��L��J
	keyo:buffer std_logic_vector(3 downto 0)	--��L��X
	);	 
end KTM626;

-- -----------------------------------------------------
architecture Albert of KTM626 is
-- ======================= �ŧi�s�� ========================
	--UART_T1 & RS232_R2
	--UART_T1--------------------------------------------
	component RS232_T1 is
	port(clk,Reset:in std_logic;			
		--clk:25MHz
		DL:in std_logic_vector(1 downto 0);
	 	--00:5,01:6,10:7,11:8 Bit
		ParityN:in std_logic_vector(2 downto 0);
		--000:None,100:Even,101:Odd,110:Space,111:Mark
		StopN:in std_logic_vector(1 downto 0);
		--0x:1Bit,10:2Bit,11:1.5Bit
		F_Set:in std_logic_vector(2 downto 0); --�j�v�]�w
		Status_s:out std_logic_vector(1 downto 0);
		TX_W:in std_logic;
		TXData:in std_logic_vector(7 downto 0);
		TX:out std_logic);
	end component RS232_T1;
	--UART_R2--------------------------------------------
	component RS232_R2 is
	port(Clk,Reset:in std_logic;--clk:25MHz
		DL:in std_logic_vector(1 downto 0);
	 	--00:5,01:6,10:7,11:8 Bit
		ParityN:in std_logic_vector(2 downto 0);
		--0xx:None,100:Even,101:Odd,110:Space,111:Mark
		StopN:in std_logic_vector(1 downto 0);
		--0x:1Bit,10:2Bit,11:1.5Bit
		F_Set:in std_logic_vector(2 downto 0); --�j�v�]�w
		Status_s:out std_logic_vector(2 downto 0);
		Rx_R:in std_logic;
		RD:in std_logic;
		RxDs:out std_logic_vector(7 downto 0));
	end component RS232_R2;
	--�ŧiUART�`�ƻP�H��-------------------------------
	constant DL:std_logic_vector(1 downto 0):="11";
	--00:5,01:6,10:7,11:8 Bit
	constant ParityN:std_logic_vector(2 downto 0):="000";
	--0xx:None,100:Even,101:Odd,110:Space,111:Mark
	constant StopN:std_logic_vector(1 downto 0):="00";
	--0x>1Bit,10>2Bit,11>1.5Bit
	constant F_Set:std_logic_vector(2 downto 0):="101";
	--9600 BaudRate
	
	signal S_RESET_T:std_logic;		--UART�ǿ魫�m
	signal TX_W:std_logic;
	signal Status_Ts:std_logic_vector(1 downto 0);
	signal TXData:std_logic_vector(7 downto 0);
	
	signal S_RESET_R:std_logic;		--UART�������m
	signal Rx_R:std_logic;
	signal Status_Rs:std_logic_vector(2 downto 0);
	signal RxDs:std_logic_vector(7 downto 0);
	
	signal RD:std_logic;
	signal TX:std_logic;
	
	
	signal CMDn,CMDn_R:integer range 0 to 3;--UART�ǥX��,������
	--�W��PC���(4 byte)
	type pc_up_data_T is array(0 to 3) of std_logic_vector(7 downto 0);
	--�R�O
	signal pc_up_data:pc_up_data_T:=("00000000","00000000","00000000","00000000");
	
	constant hTemp:integer:=28;
	
	--DHT11�Ʀ����׷P����--------------------------------------------
	--Data format:
	--DHT11_DBo(std_logic_vector:8bit):��DHT11_RDp�����X��
	--RDp=5:chK_SUM
	--RDp=4 + 3 + 2 + 1 + 0
	--4:���(���)+3:���(�p��)+�ū�(���)+�ū�(�p��)+�P���ˬd
	--������X���(DHT11_DBoH)�ηū�(DHT11_DBoT):integer(0~255:8bit)
	component DHT11_driver is
		port(DHT11_CLK,DHT11_RESET:in std_logic;
			--DHT11_CLK:781250Hz(50MHz/2^6:1.28us:FD(5))�ާ@�t�v,���m
			DHT11_D_io:inout std_logic;			--DHT11 i/o
			DHT11_DBo:out std_logic_vector(7 downto 0);	
			--DHT11_driver ��ƿ�X
			DHT11_RDp:in integer range 0 to 7;	--���Ū������
			DHT11_tryN:in integer range 0 to 7;	--���~����մX��
			DHT11_ok,DHT11_S:buffer std_logic;
			--DHT11_driver�����@�~�X��,���~�H��
			DHT11_DBoH,DHT11_DBoT:out integer range 0 to 255);
			--������X��פηū�
	end component DHT11_driver;

	signal DHT11_CLK,DHT11_RESET:std_logic;
	--DHT11_CLK:781250Hz(50MHz/2^6:1.28us:FD(5))�ާ@�t�v,���m
	signal DHT11_DBo:std_logic_vector(7 downto 0);	--DHT11_driver ��ƿ�X
	signal DHT11_RDp:integer range 0 to 7;		--���Ū������5~0
	signal DHT11_tryN:integer range 0 to 7:=3;	--���~����մX��
	signal DHT11_ok,DHT11_S:std_logic;
	--DHT11_driver�����@�~�X��,���~�H��	
	signal DHT11_DBoH,DHT11_DBoT:integer range 0 to 255;--������X��פηū�
	
	--WS2812B��C��LED�X�ʾ�--------------
	component WS2812B_Driver is
		port(WS2812BCLK,WS2812BRESET,loadck:in std_logic;
			--�ާ@�W�v,���m,���Jck
			LEDGRBdata:in std_logic_vector(23 downto 0);
			--��m���
			reload,emitter,WS2812Bout:out std_logic);
			--�n�D���J,�o�g���A,�o�g��X 
	end component WS2812B_Driver;

	signal WS2812BCLK,WS2812BRESET,loadck,reload,emitter:std_logic;
	--�ާ@�W�v,���m,���Jck,�n�D���J,�o�g���A
	signal LEDGRBdata:std_logic_vector(23 downto 0);--��m���
	--------------------------------------------------------------------
	signal FD2:std_logic_vector(3 downto 0);
	--WS2812B_Driver���W��
	signal SpeedS,WS2812BPCK:std_logic;
	--WS2812BP�ާ@�W�v���,WS2812BP�ާ@�W�v
	signal delay:integer range 0 to 127;			--����ɶ�
	signal LED_WS2812B_N:integer range 0 to 127;	--WS2812B�Ӽƫ���
	constant NLED:integer range 0 to 127:=29;
	--WS2812B�Ӽ�:30��(0~29)
	signal LED_WS2812B_shiftN:integer range 0 to 7;	
	--WS2812B����Ӽƫ���
	signal dir_LR:std_logic_vector(15 downto 0);   	--��V����
	type LED_T is array(0 to 7) of std_logic_vector(23 downto 0);
	--�Ϲ��榡
	--�Ϲ�
	signal LED_WS2812B_T8:LED_T:=(
					"000000001111111100000000",
					"111111110000000000000000",
					"000000000000000011111111",
					"000000000000000000000000",
					"111111111111111100000000",
					"000000001111111111111111",
					"111111110000000011111111",
					"111111111111111111111111");
								
	--MG90S���A���X�ʾ�--------------
	component MG90S_Driver is
	port(MG90S_CLK,MG90S_RESET:in std_logic;
		--MG90S_Driver�X��clk(6.25MHz),reset�H��
		MG90S_dir0:in std_logic;			--��ʤ�V0
		MG90S_deg0:in integer range 0 to 90;	--��ʨ���0
		MG90S_o0:out std_logic;				--Driver��X0
		MG90S_dir1:in std_logic;			--��ʤ�V1
		MG90S_deg1:in integer range 0 to 90;	--��ʨ���1
		MG90S_o1:out std_logic);			--Driver��X1
	end component MG90S_Driver;
	signal MG90S_CLK,MG90S_RESET:std_logic;
	--MG90S_Driver�X��clk(25MHz),reset�H��
	signal MG90S_dir0,MG90S_dir1:std_logic;	--��ʤ�V
	signal MG90S_deg0,MG90S_deg1:integer range 0 to 90;
	--��ʨ���
	
	--RGB16x16 �m��ݪO-------------------
	component RGB16x16_EP3C16Q240C8 is
--	port(gckp31,SResetp99:in std_logic;	--�t���W�v,�t��reset
	port(gckp31,RGB16x16Reset:in std_logic;	--�t���W�v,�t��reset
		--DM13A
		DM13ACLKo:out std_logic;
		DM13ASDI_Ro,DM13ASDI_Go,DM13ASDI_Bo:out std_logic;
		DM13ALEo,DM13AOEo:out std_logic;
		--Scan
		Scan_DCBAo:buffer std_logic_vector(3 downto 0) );
	end component RGB16x16_EP3C16Q240C8;
	
	-- ADC ---------------------------
	component MCP3202_Driver is
	port(MCP3202_CLK_D,MCP3202_RESET:in std_logic;
		--MCP3202_Driver�X��clk,reset�H��
		MCP3202_AD0,MCP3202_AD1:buffer integer range 0 to 4095;
		--MCP3202 AD0,1 ch0,1��
		MCP3202_try_N:in integer range 0 to 3;	--���ѫ�A���զ���
		MCP3202_CH1_0:in std_logic_vector(1 downto 0);--��J�q�D
		MCP3202_SGL_DIFF:in std_logic;	--MCP3202 SGL/DIFF
		MCP3202_Do:in std_logic;		--MCP3202 do�H��
		MCP3202_Di:out std_logic;		--MCP3202 di�H��
		MCP3202_CLK,MCP3202_CS:buffer std_logic;
		--MCP3202 clk,/cs�H��
		MCP3202_ok,MCP3202_S:buffer std_logic);
		--Driver�����X�� ,�������A
	end component MCP3202_Driver;
	
	signal MCP3202_CLK_D,MCP3202_RESET:std_logic;
	--MCP3202_Driver�X��clk,reset�H��
	signal MCP3202_AD0,MCP3202_AD1:integer range 0 to 4095;
	--MCP3202 AD��
	signal MCP3202_try_N:integer range 0 to 3:=1;
	--���ѫ�A���զ���
	signal MCP3202_CH1_0:std_logic_vector(1 downto 0):="01";--ch1
	signal MCP3202_SGL_DIFF:std_logic:='1';
	--MCP3202 SGL/DIFF ��SGL
	signal MCP3202_ok,MCP3202_S:std_logic;		
	--Driver�����X�� ,�������A
	
	--timer�Ʀ����---------------------
	component timer0 is
	port(GCKP31,SResetP99,p20s1,p21s2: in std_logic;
		scan:buffer unsigned(3 downto 0);			--���˫H��
		D7data:out std_logic_vector(6 downto 0);	--��ܸ��
		D7xx_xx:out std_logic	);				--:
	end component timer0;
	
	--ROTATE_ENCODER-����s�X��------------------------
	component ROTATE_ENCODER_EP3C16Q240C8 is 
	port(gckp31,ROTATEreset:in std_logic;	--�t���W�v,�t��reset
		APi,BPi,PBi:in std_logic;
		rsw:buffer std_logic_vector(2 downto 0));--3�줸�p�ƾ�
	end component ROTATE_ENCODER_EP3C16Q240C8;
	signal ROTATEreset:std_logic;				--���m
	
	--4x4��L----------------------------------
	component KEYboard_EP3C16Q240C8 is
	port(gckp31,KEYboardreset:in std_logic;		--�t���W�v,�t��reset
		keyi:in std_logic_vector(3 downto 0);	--��L��J
		keyo:buffer std_logic_vector(3 downto 0);	--��L��X
		ksw:out std_logic_vector(2 downto 0) 	);	--0~7���
	end component KEYboard_EP3C16Q240C8;
	signal KEYboardreset:std_logic;				--���m

	----------------------------------------------------------------
	--����LCM 4bit�X�ʾ�(WG14432B5)
	component LCM_4bit_driver is
	port(LCM_CLK,LCM_RESET:in std_logic;	--�ާ@�t�v,���m
		RS,RW:in std_logic;				--�Ȧs�����,Ū�g�X�п�J
		DBi:in std_logic_vector(7 downto 0);	--LCM_4bit_driver ��ƿ�J
		DBo:out std_logic_vector(7 downto 0);	--LCM_4bit_driver ��ƿ�X
		DB_io:inout std_logic_vector(3 downto 0);	--LCM DATA BUS����
		RSo,RWo,Eo:out std_logic;		--LCM �Ȧs�����,Ū�g,�P�श��
		LCMok,LCM_S:out boolean	);		--LCM_8bit_driver����,���~�X��
	end component LCM_4bit_driver;

	signal LCM_RESET,RS,RW:std_logic;		
	--LCM_4bit_driver���m,LCM�Ȧs�����,Ū�g�X��
	signal DBi,DBo:std_logic_vector(7 downto 0);
	--LCM_4bit_driver�R�O�θ�ƿ�J�ο�X
	signal LCMok,LCM_S:boolean;			
	--LCM_4bit_driver�����@�~�X��,���~�H��

	----����LCM���O&��ƪ�榡:
	----(�`��,���O��,���O...���...........
	----�^�ƫ�LCM 4�줸�ɭ�,2�C���

	type LCM_T is array (0 to 20) of std_logic_vector(7 downto 0);
	constant LCM_IT:LCM_T:=(X"15",X"06",----���嫬LCM 4�줸�ɭ�
						"00101000","00101000","00101000",--4�줸�ɭ�
						"00000110","00001100","00000001",
						--ACC+1��ܹ��L����,��ܹ�on�L��еL�{�{,�M����ܹ�
--	X"01",X"48",X"65",X"6C",X"6C",X"6F",X"21",X"20",X"20",X"20",x"20",X"20",X"20");
--	--Hello!
	X"4B", X"54", X"4D", X"36", X"32", X"36",	--KTM626
	X"B9", X"C5",  X"A6", X"7E",  X"B5", X"D8",	--�Ŧ~��
	X"20");--�ť�

	--LCM=1:�Ĥ@�C��ܰ� LEDx16�]���O�q
	constant LCM_1:LCM_T:=(	X"15",X"01",			--�`��,���O��
						"00000001",			--�M����ܹ�
						--��1�C��ܸ��
	X"4C",X"45",X"44",X"78",X"31",X"36",X"B6",X"5D",X"B0",X"A8",X"BF",X"4F",X"A8",X"71",
	X"20",X"20",X"20",X"20");--LEDx16�]���O�q
							
	--LCM=2:�Ĥ@�C��ܰ� ����IC�θ��ﾹ����
	constant LCM_2:LCM_T:=(	X"15",X"01",			--�`��,���O��
						"00000001",			--�M����ܹ�
						--��1�C��ܸ��
	X"AD",X"B5",X"BC",X"D6",X"49",X"43",X"A4",X"CE",X"B8",X"C1", --����IC�θ��ﾹ����
	X"BB",X"EF",X"BE",X"B9",X"B4",X"FA",X"B8",X"D5");--����IC�θ��ﾹ����
	
	--LCM=3:�Ĥ@�C��ܰ� DHT11 ����״���
	signal LCM_3:LCM_T:=(	X"15",X"01",			--�`��,���O��
						"00000001",			--�M����ܹ�
						--��1�C��ܸ��
	X"44",X"48",X"54",X"31",X"31",X"20",X"B7",X"C5",X"C0",X"E3", --DHT11 ����״���
	X"AB",X"D7",X"B4",X"FA",X"B8",X"D5",X"20",X"20");--DHT11 ����״���

	--LCM=32:�ĤG�C��ܰ� �ū�  �J���  %RH
	signal LCM_32:LCM_T:=(	X"15",X"01",			--�`��,���O��
						"10010000",			--�]�ĤG�CACC��m
						--��2�C��ܸ��
	X"B7",X"C5",X"AB",X"D7",X"20",X"20",X"A2",X"4A",X"C0",X"E3",--�ū�  �J���  %RH
	X"AB",X"D7",X"20",X"20",X"25",X"52",X"48",X"20");--�ū�  �J���  %RH
	
	--LCM=4:�Ĥ@�C��ܰ� WS2812B RGB ����
	constant LCM_4:LCM_T:=(	X"15",X"01",			--�`��,���O��
						"00000001",			--�M����ܹ�
						--��1�C��ܸ��
	X"57",X"53",X"32",X"38",X"31",X"32",X"42",X"20",X"52",X"47", --WS2812B RGB ���� 
	X"42",X"20",X"B4",X"FA",X"B8",X"D5",X"20",X"20");--WS2812B RGB ���� 
							
	--LCM=5:�Ĥ@�C��ܰ� �����u���� 
	constant LCM_5:LCM_T:=(	X"15",X"01",			--�`��,���O��
						"00000001",			--�M����ܹ�
						--��1�C��ܸ��
	X"BE",X"F7",X"B1",X"F1",X"C1",X"75",X"B4",X"FA",X"B8",X"D5",--�����u����
	X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20");--�����u���� 
							
	--LCM=6:�Ĥ@�C��ܰ� RGB16x16�q
	constant LCM_6:LCM_T:=(	X"15",X"01",			--�`��,���O��
						"00000001",			--�M����ܹ�
						--��1�C��ܸ��
	X"52",X"47",X"42",X"31",X"36",X"78",X"31",X"36",X"A8",X"71",--RGB16x16�q
	X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20");--RGB16x16�q
							
	--LCM=7:�Ĥ@�C��ܰ� LM35 �ū״���
	constant LCM_7:LCM_T:=(	X"15",X"01",			--�`��,���O��
						"00000001",			--�M����ܹ�
						--��1�C��ܸ��
	X"4C",X"4D",X"33",X"35",X"B7",X"C5",X"AB",X"D7",X"B4",X"FA",--LM35 �ū״���
	X"B8",X"D5",X"20",X"20",X"20",X"20",X"20",X"20");--LM35 �ū״���
							
	--LCM=72:�ĤG�C��ܰ� �ū�xxx.x�J
	signal LCM_72:LCM_T:=(	X"15",X"01",			--�`��,���O��
						"10010000",			--�]�ĤG�CACC��m
						--��2�C��ܸ��
	X"B7",X"C5",X"AB",X"D7",X"20",X"20",X"20",X"2E",X"20",X"20",--�ū�xxx.x�J
	X"A2",X"4A",X"20",X"20",X"20",X"20",X"20",X"20");--�ū�xxx.x�J
							
	signal LCM_com_data,LCM_com_data2:LCM_T;
	signal LCM_INI:integer range 0 to 31;
	signal LCMP_RESET,LN,LCMPok:std_logic;
	signal LCM,LCMx:integer range 0 to 7;
	
----- �ŧi��L�H�� ---------------
	signal FD:std_logic_vector(30 downto 0);	--���W��
	signal times:integer range 0 to 2047;		--�p�ɾ�
	signal S0S,S1S,S2S,M0S,M1S,M2S:std_logic_vector(2 downto 0);
	--S0,S1,S2,M0,M1,M2���u��
	signal MMx,MM,PCswx,rsw,ksw:std_logic_vector(2 downto 0);
	signal LED_LR_dir,SW_CLK,sound1on,LCD_refresh,WS2812BPReset:std_logic;
	signal MG90S_sch,MG90S_s,RGB16x16Reset:std_logic;
	signal autoMM:std_logic_vector(2 downto 0);
	signal lm35T:integer range 0 to 1550;
begin
---- �s�� RS232�s�� -------------------
--RS232�ǰe�Ҳ�
U1: RS232_T1 
	port map(FD(0),S_RESET_T,DL,ParityN,StopN,F_Set,Status_Ts,TX_W,TXData,TX);
--RS232�����Ҳ�	
U2: RS232_R2
	port map(FD(0),S_RESET_R,DL,ParityN,StopN,F_Set,Status_Rs,Rx_R,RD,RxDs);			

---- �s�� DHT11�s�� -------------------
DHT11_CLK<=FD(5);	--DHT11_CLK:781250Hz(50MHz/2^6:1.28us:FD(5))�ާ@�t�v
U3: DHT11_driver
	port map(	DHT11_CLK,DHT11_RESET,
--DHT11_CLK:781250Hz(50MHz/2^6:1.28us:FD(5))�ާ@�t�v,���m
			DHT11_D_io,		--DHT11 i/o
			DHT11_DBo,		--DHT11_driver ��ƿ�X
			DHT11_RDp,		--���Ū������
			DHT11_tryN,		--���~����մX��
			DHT11_ok,DHT11_S,DHT11_DBoH,DHT11_DBoT);	
			--DHT11_driver�����@�~�X��,���~�H��,������X��פηū�	
---- �s�� LCM�s�� -------------------
LCMset: LCM_4bit_driver
	port map(FD(7),LCM_RESET,RS,RW,DBi,DBo,DB_io,RSo,RWo,Eo,LCMok,LCM_S);	

---- �s�� WS2812B�s�� -------------------
WS2812BN: WS2812B_Driver
	port map(	WS2812BCLK,WS2812BRESET,loadck,LEDGRBdata,
			reload,emitter,WS2812Bout);
		  	WS2812BRESET<=SResetP99;	--�t��reset

---- �s�� MG90S�s�� -------------------
MG90S: MG90S_Driver
 	port map(	FD(2),MG90S_RESET,--MG90S_Driver�X��clk(6.25MHz),reset�H��
			MG90S_dir0,	--��ʤ�V0
			MG90S_deg0,	--��ʨ���0
			MG90S_o0,	--Driver��X0
			MG90S_dir1,	--��ʤ�V1
			MG90S_deg1,	--��ʨ���1
			MG90S_o1);	--Driver��X1
						  
---- �s�� RGB16x16�s�� -------------------
RGB16x16:RGB16x16_EP3C16Q240C8 
	port map(	gckp31,RGB16x16Reset,	--�t���W�v,RGB16x16Reset
			--DM13A
			DM13ACLKo,
			DM13ASDI_Ro,DM13ASDI_Go,DM13ASDI_Bo,
			DM13ALEo,DM13AOEo,
			--Scan
			Scan_DCBAo);

---- �s�� MCP3202�s�� -------------------
U4: MCP3202_Driver
	port map(	FD(4),MCP3202_RESET,	--MCP3202_Driver�X��clk,reset�H��
			MCP3202_AD0,MCP3202_AD1,--MCP3202 AD��
			MCP3202_try_N,			--���ѫ�A���զ���
			MCP3202_CH1_0,			--��J�q�D
			MCP3202_SGL_DIFF,		--SGL/DIFF
			MCP3202_Do,			--MCP3202 do�H��
			MCP3202_Di,			--MCP3202 di�H��
			MCP3202_CLK,MCP3202_CS,	--MCP3202 clk,/cs�H�� 
			MCP3202_ok,MCP3202_S);	--Driver�����X�� ,�������A

---- �s�� ���� �s�� -------------------
U5:timer0 port map(	GCKP31,SResetP99,PB7,PB8,
				scan, D7data,		--���˫H���B��ܸ��
		  		D7xx_xx);			--:�{��
				   
---- �s�� ����s�X�� �s�� -------------------
U6:ROTATE_ENCODER_EP3C16Q240C8 
	port map(	gckp31,ROTATEreset,		--�t���W�v,�t��reset
			APi,BPi,PBi,
			rsw	);
	
---- �s�� 4x4��L �s�� -------------------
U7:KEYboard_EP3C16Q240C8
	port map(	gckp31,KEYboardreset,--�t���W�v,�t��reset
			keyi, keyo,		--��L��J�B��L��X
			ksw);			--0~7���

--------------------------------------------------------------------------
-- �z�Luart�W�ǷūסB��׸��
TXData<=pc_up_data(CMDn-1);
pc_up_data(1)<=	conv_std_logic_vector(DHT11_DBoT,8) when MM="011" else
 				conv_std_logic_vector(MCP3202_AD1/256,8);
				--�W��PC��� DHT11 �ū� or LM35 ADC
pc_up_data(0)<=	conv_std_logic_vector(DHT11_DBoH,8) when MM="011" else
 				conv_std_logic_vector(MCP3202_AD1 mod 256,8);
				--�W��PC��� DHT11 ��� or LM35 ADC

------------------------------------------------------
UART_command_Main:process(FD(17))
begin
	if SResetP99='0' then		--�t�έ��m
		Rx_R<='0';			--����Ū���H��
		TX_W<='0';			--������Ƹ��J�H��
		S_RESET_T<='0';		--����UART�ǰe
		S_RESET_R<='0';		--����UART����
		CMDn<=0;				--�W��0byte
		CMDn_R<=1;			--�����ƶq(1byte)
		PCswx<="000";
	elsif (Rx_R='1' and Status_Rs(2)='0') then	--UART�����Y�ɳB�z
		Rx_R<='0';						--�Y�ɨ���Ū���H��
	elsif rising_edge(FD(17)) then
		S_RESET_T<='1';				--�}��UART�ǰe
		S_RESET_R<='1';				--�}��UART����
		if CMDn>0 and S_RESET_T='1' then	--�W��
			if Status_Ts(1)='0' then	--�ǰe�w�İϤw��
				if TX_W='1' then
					TX_W<='0';		--�����ǰe��Ƹ��J�ɯ�
					CMDn<=CMDn-1;		--���Ы��V�U�@�����
				else
					TX_W<='1';		--�ǰe��Ƹ��J�ɯ�
				end if;
			end if;
		-----------------------
		--�w������UART�R�O
		elsif Status_Rs(2)='1' then		--�w������UART�R�O
			Rx_R<='1';				--Ū���H��
			--PC�R�O�ѪR-------------------
			PCswx<=RxDs(2 downto 0);	--����UART�R�O
		end if;
		
		if 	(MM="011" and LCD_refresh='1' and DHT11_ok='1') or
	 		(MM="111" and LCD_refresh='1' and MCP3202_ok='1') then CMDn<=2;	
			--�W��2byte(�W�� DHT11 �����)
		end if;
	end if;
end process UART_command_Main;

--on(0)=USB, off(1)=BT(����)
RD <= USB_TX when dip15P57='0' else BT_TX;
USB_RX <= TX when dip15P57='0' else 'Z';
BT_RX <= TX when dip15P57='1' else 'Z';	

--�\��۰ʮi�ܤ���-----------------------------------------------------------------------------------
autoswitch:process(FD(30))
begin
	if S0S(2)='0' then
		autoMM<="000";		--�q��1�ӥ\��}�l
	elsif rising_edge(FD(30)) then	
		autoMM<=autoMM+1; 	--�U�@�ӥ\��
	end if;
end process autoswitch;
------------------------------------
MMx<=autoMM when S0S(2)='1' else 
M2S(2)& M1S(2)& M0S(2)	when S1S(2)='0' and S2S(2)='0' else 
	rsw 				when S1S(2)='0' and S2S(2)='1' else 
	ksw					when S1S(2)='1' and S2S(2)='0' else
 	PCswx;--����R�O�ӷ�:�����}����PC 

KTM626_Main:process(FD(17))
begin
	if SResetP99='0' then	--�t�έ��m
		MM<=not MMx;		--���������}���������������}�����A
		led16<=(others=>'1');--����16��LED
		LCMP_RESET<='0';
		LCM<=0;
		sound1on<='0';
		sound2<='0';
		DHT11_RESET<='0';
		WS2812BPReset<='0';
		MG90S_RESET<='0';
		RGB16x16Reset<='0';
		MCP3202_RESET<='0';
		ROTATEreset<='0';
		KEYboardreset<='0';
	elsif rising_edge(FD(17)) then
		LCMP_RESET<='1';
		ROTATEreset<='1';
		KEYboardreset<='1';
		if LCMPok='1' then
			if MM/=MMx then	-- �����i�ܼҦ�
			--��������}����������������}�����A�δ��յ{�ǰ���(����S1)
				MM<=MMx;			
				--���������}�������������}�����A
				DHT11_RESET<='0';		--DHT11_driver����X��
				led16<=(others=>'1');	--����16��LED
				sound1on<='0'; 			--�������ﾹ1
				sound2<='0'; 			--�������ﾹ2(����IC)
				WS2812BPReset<='1'; 	--��C��LED����X��
				MG90S_RESET<='0'; 		--���A������X��
				RGB16x16Reset<='0'; 	--RGB�ݪO����X��
				MCP3202_RESET<='0'; 	--ADC����X��
				case MMx is			--�ھګ����}�����A
					when "001" =>	--001:LED16�q
						LED_LR_dir<='0';--�]�wLED��V
						led16<=(others=>'0');--����16��LED
						times<=10; 	--�]�w����LED16�q����
						LCM<=1; 		--LCD���
					when "010" =>	--010:���ﾹ��X
						LCM<=2; 		--LCD���
						times<=200; 	--�]�w���榸��
					when "011" =>	--011:DHT11 ����״���
						LCM<=3; 		--LCD���
						times<=800; 	--�]�w���榸��
					when "100" =>	--100:WS2812B��C��LED�q
						WS2812BPReset<='0';
						LCM<=4; 		--LCD���
					when "101" =>	--101:MG90S���A���q
						LCM<=5; 		--LCD���
						MG90S_dir0<='0';--�]�w�Ĥ@�x���A������ʤ�V0
						MG90S_deg0<=0;	--�]�w�Ĥ@�x���A������ʨ���0
						MG90S_dir1<='0';--�]�w�ĤG�x���A������ʤ�V1
						MG90S_deg1<=0;	--�]�w�ĤG�x���A������ʨ���1
						times<=10; 	--�]�w���榸��
						MG90S_s<='0'; 	--�]�w�Ĥ@�x���A���}�l����
						MG90S_sch<='0';--�]�w���楿��
					when "110" =>	--110: RGB16x16�m��ݪO�q
						LCM<=6; 		--LCD���
					when "111" =>	--111:LM35����ū״���
						LCM<=7; 		--LCD���
						times<=500; 	--�]�w���榸��
					when others =>	--000:����
					
						LED_LR_dir<='0';--�]�wLED��V
						led16<=(others=>'0');--����16��LED
						times<=10; 	--�]�w����LED16�q����

						WS2812BPReset<='0';

						MG90S_dir0<='0';--�]�w�Ĥ@�x���A������ʤ�V0
						MG90S_deg0<=0;	--�]�w�Ĥ@�x���A������ʨ���0
						MG90S_dir1<='0';--�]�w�ĤG�x���A������ʤ�V1
						MG90S_deg1<=0;	--�]�w�ĤG�x���A������ʨ���1
						times<=10; 	--�]�w���榸��
						MG90S_s<='0'; 	--�]�w�Ĥ@�x���A���}�l����
						MG90S_sch<='0';--�]�w���楿��
					
						LCM<=0; 		--LCD���

				end case;
			else		-- ����i�ܼҦ�
				times<=times-1;
				case MMx is
				
				
					---000-----------------------------------
					--	MG90S_dir0=0�B	MG90S_deg0=0
					--	MG90S_dir1=0�B	MG90S_deg1=0
					--	times=10�BMG90S_s=0(�Ĥ@�x)�BMG90S_sch=0(����)
					--	LCM<=5 
					when "000" =>	--101:MG90S���A������
						
						if times=0 then
							times<=10;
							if LED_LR_dir='1' then
								led16<=led16(14 downto 0) & not led16(15);	
								--16bit����:�j�ͧުk
								LED_LR_dir<=led16(15) or not led16(14);
							else
								led16<=not led16(0) & led16(15 downto 1);	
								--16bit�k��:�j�ͧުk
								LED_LR_dir<=led16(1) and not led16(0);	
							end if;
						end if;
						
						if dip16P56='0' then
							sound2<='1'; ---����IC�s��
						else
							sound2<='0'; ---����IC���s��
						end if;

						RGB16x16Reset<='1'; --���ҬݪO

						WS2812BPReset<='1';
					
						MG90S_RESET<='1';
						if times=0 then
							times<=3;
							if MG90S_s='0' then
							--�ާ@�Ĥ@�x���A��
								if MG90S_sch='0' then
								--����
									MG90S_deg0<=MG90S_deg0+1;
									if MG90S_deg0=90 then
										MG90S_deg0<=89;
										MG90S_sch<='1';
									end if;
								else
								--����
									MG90S_deg0<=MG90S_deg0-1;
									if MG90S_deg0=0 then
										MG90S_deg0<=0;
										MG90S_dir0<=not MG90S_dir0;
										MG90S_sch<='0';
										MG90S_s<=MG90S_dir0;
									end if;
								end if;
							else
							--�ާ@�ĤG�x���A��
								if MG90S_sch='0' then
								--����
									MG90S_deg1<=MG90S_deg1+1;
									if MG90S_deg1=90 then
										MG90S_deg1<=89;
										MG90S_sch<='1';
									end if;
								else
								--����
									MG90S_deg1<=MG90S_deg1-1;
									if MG90S_deg1=0 then
										MG90S_deg1<=0;
										MG90S_dir1<=not MG90S_dir1;
										MG90S_sch<='0';
										MG90S_s<=not MG90S_dir1;
									end if;
								end if;
							end if;											
						end if;
				
				
					---001-----------------------------------
					--	LED_LR_dir=0�Bled16=0�Btimes=10 
					--	LCM=1 
					when "001" =>	--LED16  --�Ӧ^:�j�ͧުk
						if times=0 then
							times<=10;
							if LED_LR_dir='1' then
								led16<=led16(14 downto 0) & not led16(15);	
								--16bit����:�j�ͧުk
								LED_LR_dir<=led16(15) or not led16(14);
							else
								led16<=not led16(0) & led16(15 downto 1);	
								--16bit�k��:�j�ͧުk
								LED_LR_dir<=led16(1) and not led16(0);	
							end if;
						end if;
	
					---010-----------------------------------
					--	times=200�BLCM=2
					when "010" =>	--���ﾹ��X
						---sound1�Psound2���O�ߪi�����ﾹ(���A�ʧ@)
						---sound2�ѭ���IC�X��
						--if times=40 then	---�ͤ@�n
						--	sound1on<='1';
						--end if;
						--if times=0 then
						--	sound1on<='0';
						--	times<=200;
						--end if;
						sound2<='1'; ---����IC
						
					---011-----------------------------------
					--	times=800�BLCM=3
					when "011" =>	--DHT11 ����״���
					
						if dip16P56='0' then
							sound2<='1'; ---����IC�s��
						else
							sound2<='0'; ---����IC���s��
						end if;
					
					
						if DHT11_RESET='0' then	--DHT11_driver�|���Ұ�
							DHT11_RESET<='1';	--DHT11���Ū��
							LCD_refresh<='1'; 	--��sLCD�X�г]�w��1
						elsif DHT11_ok='1' then	--DHT11Ū������
							if LCD_refresh='1' then--��sLCD�W�������
								LCMP_RESET<='0'; --����LCD 
								LCD_refresh<='0';--��sLCD�X�г]�w��0
								times<=800;
							elsif times=0 then
								DHT11_RESET<='0';	--DHT11�ǳƭ��sŪ�����
							elsif DHT11_S='1' then	--���Ū������
								null;			--�ƻ򳣧O��(����)
							elsif DHT11_DBoT>hTemp then--�ū׶W�LhTemp��
								sound1on<='1'; 	--�ͤ@�n
							else
								sound1on<='0';
							end if;
						end if;
	
					---100-----------------------------------
					--	WS2812BPReset=0
					--	LCM=4
					when "100"  =>	--WS2812B��C��LED�q
						WS2812BPReset<='1';

						if dip16P56='0' then
							sound2<='1'; ---����IC�s��
						else
							sound2<='0'; ---����IC���s��
						end if;


					---101-----------------------------------
					--	MG90S_dir0=0�B	MG90S_deg0=0
					--	MG90S_dir1=0�B	MG90S_deg1=0
					--	times=10�BMG90S_s=0(�Ĥ@�x)�BMG90S_sch=0(����)
					--	LCM<=5 
					when "101" =>	--101:MG90S���A������
						MG90S_RESET<='1';
						if times=0 then
							times<=3;
							if MG90S_s='0' then
							--�ާ@�Ĥ@�x���A��
								if MG90S_sch='0' then
								--����
									MG90S_deg0<=MG90S_deg0+1;
									if MG90S_deg0=90 then
										MG90S_deg0<=89;
										MG90S_sch<='1';
									end if;
								else
								--����
									MG90S_deg0<=MG90S_deg0-1;
									if MG90S_deg0=0 then
										MG90S_deg0<=0;
										MG90S_dir0<=not MG90S_dir0;
										MG90S_sch<='0';
										MG90S_s<=MG90S_dir0;
									end if;
								end if;
							else
							--�ާ@�ĤG�x���A��
								if MG90S_sch='0' then
								--����
									MG90S_deg1<=MG90S_deg1+1;
									if MG90S_deg1=90 then
										MG90S_deg1<=89;
										MG90S_sch<='1';
									end if;
								else
								--����
									MG90S_deg1<=MG90S_deg1-1;
									if MG90S_deg1=0 then
										MG90S_deg1<=0;
										MG90S_dir1<=not MG90S_dir1;
										MG90S_sch<='0';
										MG90S_s<=not MG90S_dir1;
									end if;
								end if;
							end if;											
						end if;
	
					---110-----------------------------------
					--	LCM=6
					when "110" =>	--RGB16x16 test
						RGB16x16Reset<='1'; --���ҬݪO
						
					---111-----------------------------------
					--	times=500�BLCM=7
					when "111" =>	--LM35����ū׷P��
						if MCP3202_RESET='0' then	--LM35_driver�|���Ұ�
							MCP3202_RESET<='1';		--LM35���Ū��
							LCD_refresh<='1';
						elsif MCP3202_ok='1' then	--LM35Ū������
							if LCD_refresh='1' then
								LCMP_RESET<='0';
								LCD_refresh<='0';
								times<=500;
							elsif times=0 then		--�ɶ���
								MCP3202_RESET<='0';	--LM35�ǳƭ��sŪ�����
							elsif MCP3202_S='1' then--���Ū������
								null;			--���򳣤���(����)
							end if;
						end if;
						
						if dip16P56='0' then
							sound2<='1'; ---����IC�s��
						else
							sound2<='0'; ---����IC���s��
						end if;
						
						
					when others =>--���򳣤���(����)
						null;
				end case;
			end if;
		end if;
	end if;
end process KTM626_Main;

--- ���n ---------------------------------------------------
sound1<=FD(20)and FD(16)and FD(11)and sound1on when MM="010" else FD(22)and FD(16) and sound1on;
------------------------------------------------------------
--DHT11 LCM���
LCM_32(16)<="0011" & conv_std_logic_vector(DHT11_DBoH mod 10,4);		
-- �^����פ��Ӧ��(ASCII)
LCM_32(15)<="0011" & conv_std_logic_vector((DHT11_DBoH/10)mod 10,4);	
-- �^����פ��Q���(ASCII)
LCM_32(8)<="0011" & conv_std_logic_vector(DHT11_DBoT mod 10,4);		
-- �^���ūפ��Ӧ��(ASCII)
LCM_32(7)<="0011" & conv_std_logic_vector((DHT11_DBoT/10)mod 10,4);		
-- �^���ūפ��Q���(ASCII)

--LM35 LCM���
LM35T<=MCP3202_AD1*122/100;	--5/10mv=500/4095*1000=122*MCP3202_AD1/100 xxx.x
-- MCP3202��12bit ADC(0~4095)�A�q���d��0~5V
--�C��MCP3202���5/4095 V�A��5/4095*1000 mV=1.22mV
-- LM35�C�@�ק���10mV�A�Y10m/1.22�Ө��=10/1.22�Ө��
--�Y�n�NMCP3202�ഫ�᪺�ȡA�٭쬰�ūץ������H�o�ӭ�
-------------------------------------------
--MCP3202�ഫ�᪺�Ȭ�MCP3202_ADI
--�h�ū׬�MCP3202_ADI/(10/1.22)��MCP3202_ADI*0.122
--�Y�n�H�p�Ƥ@���ܡA�h��MCP3202_ADI*1.22�A��MCP3202_ADI*122/100
--------------------------------------------
LCM_72(7)<=X"20" when LM35T<1000 else "0011" & conv_std_logic_vector(LM35T/1000,4);		
-- �^���ʦ��(ASCII)
LCM_72(8)<=X"20" when LM35T<100 else "0011" & conv_std_logic_vector((LM35T/100)mod 10,4);	
-- �^���Q���(ASCII)
LCM_72(9)<="0011" & conv_std_logic_vector((LM35T/10)mod 10,4);							
-- �^���Ӧ��(ASCII)
LCM_72(10)<=X"2E";										
--.�p���I(ASCII)
LCM_72(11)<="0011" & conv_std_logic_vector(LM35T mod 10,4);	
-- �^���p��1��(ASCII)

--��m��� ----------------------------------------
LEDGRBdata<=LED_WS2812B_T8((LED_WS2812B_N+LED_WS2812B_shiftN) mod 8) 
	when MMx="100" or MMx="000" else (others=>'0');

--WS2812BP�ާ@�W�v���
WS2812BPCK<=FD(8) when SpeedS='0' else FD(17);
--- SpeedS=0�ֳt(97.7KHz)�BSpeedS=1�C�t(191Hz)
WS2812BP:process(WS2812BPCK)
begin
	if WS2812BPReset='0' then	--���m
		LED_WS2812B_N<=0;		--�q�Y�}�l
		LED_WS2812B_shiftN<=0;	--����0
		dir_LR<=(others=>'0'); 	--15..0
		loadck<='0';
		SpeedS<='0';			--�[�־ާ@�t�v
	elsif rising_edge(WS2812BPCK) then
		if loadck='0' then		--���ݸ��J
			loadck<=reload;
		elsif LED_WS2812B_N=NLED then	--NLED��WS2812B���ƶq
			SpeedS<='1';				--��C�ާ@�t�v
			if emitter='0' then			--�w����o�g
				if delay/=0 then		--�I�G�ɶ�&�ܤƳt�v
					delay<=delay-1;	--�ɶ�����
				else
					loadck<='0';		--reemitter
					LED_WS2812B_N<=0;	--�q�Y�}�l
					dir_LR<=dir_LR+1;	--��V����
					if dir_LR(7)='1' then
					--��V����C256��WS2812BPCK�����@����V����
						LED_WS2812B_shiftN<=LED_WS2812B_shiftN+1;--���컼�W
					else
						LED_WS2812B_shiftN<=LED_WS2812B_shiftN-1;--���컼��
					end if;
					SpeedS<='0';	--�[�־ާ@�t�v
				end if;
			end if;
		else
			loadck<='0';
			LED_WS2812B_N<=LED_WS2812B_N+1;	--�վ��X��m
			delay<=20;--40;
		end if;
	end if;
end process WS2812BP;

-----------------------------------------------------
--����LCM��ܾ�
--���O&��ƪ�榡: 
--(�`��,���O��,���O...���..........
LCM_P:process(FD(0))
	variable SW:Boolean;				--�R�O�θ�ƳƧ��X��
begin
	if LCM/=LCMx or LCMP_RESET='0' then	--LCM��s���
		LCMx<=LCM;
		LCM_RESET<='0';				--LCM���m
		LCM_INI<=2;					--�R�O�θ�Ư��޳]���_�I
		LN<='0';						--�]�w��X1�C
		case LCM is
			when 0=>
				LCM_com_data<=LCM_IT;	--LCM��l�ƿ�X�Ĥ@�C���Hello!
			when 1=>
				LCM_com_data<=LCM_1;	--��X�Ĥ@�C���
			when 2=>
				LCM_com_data<=LCM_2;	--��X�Ĥ@�C���
			when 3=>
				LCM_com_data<=LCM_3;	--��X�Ĥ@�C���
				LCM_com_data2<=LCM_32;	--��X�ĤG�C���
				LN<='1';				--�]�w��X2�C
			when 4=>
				LCM_com_data<=LCM_4;	--��X�Ĥ@�C���
			when 5=>
				LCM_com_data<=LCM_5;	--��X�Ĥ@�C���
			when 6=>
				LCM_com_data<=LCM_6;	--��X�Ĥ@�C���
			when 7=>
				LCM_com_data<=LCM_7;	--��X�Ĥ@�C���
				LCM_com_data2<=LCM_72;	--��X�ĤG�C���
				LN<='1';				--�]�w��X2�C
			when others =>
				LCM_com_data<=LCM_IT;	--��X�Ĥ@�C���
		end case;
		LCMPok<='0';
		SW:=False;					--�R�O�θ�ƳƧ��X��
	elsif rising_edge(FD(0)) then		
		if SW then					--�R�O�θ�ƳƧ���
			LCM_RESET<='1';			--�Ұ�LCM_4bit_driver
			SW:=False;				--���m�X��
		elsif LCM_RESET='1' then		--LCM_4bit_driver�Ұʤ�
			if LCMok then				--����LCM_4bit_driver�����ǰe
				LCM_RESET<='0';		--������LCM���m
			end if;
		elsif LCM_INI<LCM_com_data(0) then	--�R�O�θ�Ʃ|���ǧ�
			if LCM_INI<=(LCM_com_data(1)+1) then--��R�O�θ�ƼȦs��
				RS<='0';	--Instruction reg
			else
				RS<='1';	--Data reg
			end if;
			RW<='0';		--LCM�g�J�ާ@
			DBi<=LCM_com_data(LCM_INI);	--���J�R�O�θ��
			LCM_INI<=LCM_INI+1;			--�R�O�θ�Ư��ޫ���U�@��
			SW:=True;					--�R�O�θ�Ƥw�Ƨ�
		else
			if LN='1' then
				LN<='0';
				LCM_INI<=2;			--�R�O�θ�Ư��޳]���_�I
				LCM_com_data<=LCM_com_data2;--LCM��X�ĤG�C���
			else
				LCMPok<='1';			--���槹��
			end if;
		end if;
	end if;
end process LCM_P;	

-----------------------------------------
SW_CLK<=FD(19);	--���u���ާ@�t�v
process(SW_CLK)	--���u��
begin
	
	--S0���u��
	if S0='0' then
		S0S<="000";
	elsif rising_edge(SW_CLK) then
		S0S<=S0S+ not S0S(2);
	end if;
	
	--S1���u��
	if S1='0' then
		S1S<="000";
	elsif rising_edge(SW_CLK) then
		S1S<=S1S+ not S1S(2);
	end if;
	
	--S2���u��
	if S2='0' then
		S2S<="000";
	elsif rising_edge(SW_CLK) then
		S2S<=S2S+ not S2S(2);
	end if;

	--M0���u��
	if M0='0' then
		M0S<="000";
	elsif rising_edge(SW_CLK) then
		M0S<=M0S+ not M0S(2);
	end if;

	--M1���u��
	if M1='0' then
		M1S<="000";
	elsif rising_edge(SW_CLK) then
		M1S<=M1S+ not M1S(2);
	end if;
	
	--M2���u��
	if M2='0' then
		M2S<="000";
	elsif rising_edge(SW_CLK) then
		M2S<=M2S+ not M2S(2);
	end if;
	
end process;

-- ���W��----------------------------------------
Freq_Div:process(GCKP31)
begin
	if SResetP99='0' then			--�t��reset
		FD<=(others=>'0');
		FD2<=(others=>'0');
		WS2812BCLK<='0';			--WS2812BN�X���W�v
	elsif rising_edge(GCKP31) then	--50MHz
		FD<=FD+1;
		if FD2=9 then				--7~12
			FD2<=(others=>'0');
			WS2812BCLK<=not WS2812BCLK;--50MHz/20=2.5MHz T.=. 0.4us
		else
			FD2<=FD2+1;
		end if;
	end if;
end process Freq_Div;
-- ----------------------------------------------
end Albert;

